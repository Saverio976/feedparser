module xmlreplacement

pub const xml_replacement = map{
	'&#198;':                            'Æ'
	'&AElig;':                           'Æ'
	'&#38;':                             '&'
	'&AMP;':                             '&'
	'&#193;':                            'Á'
	'&Aacute;':                          'Á'
	'&Abreve;':                          'Ă'
	'&#258;':                            'Ă'
	'&#194;':                            'Â'
	'&Acirc;':                           'Â'
	'&Acy;':                             'А'
	'&#1040;':                           'А'
	'&Afr;':                             '𝔄'
	'&#120068;':                         '𝔄'
	'&#192;':                            'À'
	'&Agrave;':                          'À'
	'&Alpha;':                           'Α'
	'&#913;':                            'Α'
	'&Amacr;':                           'Ā'
	'&#256;':                            'Ā'
	'&And;':                             '⩓'
	'&#10835;':                          '⩓'
	'&Aogon;':                           'Ą'
	'&#260;':                            'Ą'
	'&Aopf;':                            '𝔸'
	'&#120120;':                         '𝔸'
	'&ApplyFunction;':                   '⁡'
	'&#8289;':                           '⁡'
	'&#197;':                            'Å'
	'&Aring;':                           'Å'
	'&Ascr;':                            '𝒜'
	'&#119964;':                         '𝒜'
	'&Assign;':                          '≔'
	'&#8788;':                           '≔'
	'&#195;':                            'Ã'
	'&Atilde;':                          'Ã'
	'&#196;':                            'Ä'
	'&Auml;':                            'Ä'
	'&Backslash;':                       '∖'
	'&#8726;':                           '∖'
	'&Barv;':                            '⫧'
	'&#10983;':                          '⫧'
	'&Barwed;':                          '⌆'
	'&#8966;':                           '⌆'
	'&Bcy;':                             'Б'
	'&#1041;':                           'Б'
	'&Because;':                         '∵'
	'&#8757;':                           '∵'
	'&Bernoullis;':                      'ℬ'
	'&#8492;':                           'ℬ'
	'&Beta;':                            'Β'
	'&#914;':                            'Β'
	'&Bfr;':                             '𝔅'
	'&#120069;':                         '𝔅'
	'&Bopf;':                            '𝔹'
	'&#120121;':                         '𝔹'
	'&Breve;':                           '˘'
	'&#728;':                            '˘'
	'&Bscr;':                            'ℬ'
	'&Bumpeq;':                          '≎'
	'&#8782;':                           '≎'
	'&CHcy;':                            'Ч'
	'&#1063;':                           'Ч'
	'&#169;':                            '©'
	'&COPY;':                            '©'
	'&Cacute;':                          'Ć'
	'&#262;':                            'Ć'
	'&Cap;':                             '⋒'
	'&#8914;':                           '⋒'
	'&CapitalDifferentialD;':            'ⅅ'
	'&#8517;':                           'ⅅ'
	'&Cayleys;':                         'ℭ'
	'&#8493;':                           'ℭ'
	'&Ccaron;':                          'Č'
	'&#268;':                            'Č'
	'&#199;':                            'Ç'
	'&Ccedil;':                          'Ç'
	'&Ccirc;':                           'Ĉ'
	'&#264;':                            'Ĉ'
	'&Cconint;':                         '∰'
	'&#8752;':                           '∰'
	'&Cdot;':                            'Ċ'
	'&#266;':                            'Ċ'
	'&Cedilla;':                         '¸'
	'&#184;':                            '¸'
	'&CenterDot;':                       '·'
	'&#183;':                            '·'
	'&Cfr;':                             'ℭ'
	'&Chi;':                             'Χ'
	'&#935;':                            'Χ'
	'&CircleDot;':                       '⊙'
	'&#8857;':                           '⊙'
	'&CircleMinus;':                     '⊖'
	'&#8854;':                           '⊖'
	'&CirclePlus;':                      '⊕'
	'&#8853;':                           '⊕'
	'&CircleTimes;':                     '⊗'
	'&#8855;':                           '⊗'
	'&ClockwiseContourIntegral;':        '∲'
	'&#8754;':                           '∲'
	'&CloseCurlyDoubleQuote;':           '”'
	'&#8221;':                           '”'
	'&CloseCurlyQuote;':                 '’'
	'&#8217;':                           '’'
	'&Colon;':                           '∷'
	'&#8759;':                           '∷'
	'&Colone;':                          '⩴'
	'&#10868;':                          '⩴'
	'&Congruent;':                       '≡'
	'&#8801;':                           '≡'
	'&Conint;':                          '∯'
	'&#8751;':                           '∯'
	'&ContourIntegral;':                 '∮'
	'&#8750;':                           '∮'
	'&Copf;':                            'ℂ'
	'&#8450;':                           'ℂ'
	'&Coproduct;':                       '∐'
	'&#8720;':                           '∐'
	'&CounterClockwiseContourIntegral;': '∳'
	'&#8755;':                           '∳'
	'&Cross;':                           '⨯'
	'&#10799;':                          '⨯'
	'&Cscr;':                            '𝒞'
	'&#119966;':                         '𝒞'
	'&Cup;':                             '⋓'
	'&#8915;':                           '⋓'
	'&CupCap;':                          '≍'
	'&#8781;':                           '≍'
	'&DD;':                              'ⅅ'
	'&DDotrahd;':                        '⤑'
	'&#10513;':                          '⤑'
	'&DJcy;':                            'Ђ'
	'&#1026;':                           'Ђ'
	'&DScy;':                            'Ѕ'
	'&#1029;':                           'Ѕ'
	'&DZcy;':                            'Џ'
	'&#1039;':                           'Џ'
	'&Dagger;':                          '‡'
	'&#8225;':                           '‡'
	'&Darr;':                            '↡'
	'&#8609;':                           '↡'
	'&Dashv;':                           '⫤'
	'&#10980;':                          '⫤'
	'&Dcaron;':                          'Ď'
	'&#270;':                            'Ď'
	'&Dcy;':                             'Д'
	'&#1044;':                           'Д'
	'&Del;':                             '∇'
	'&#8711;':                           '∇'
	'&Delta;':                           'Δ'
	'&#916;':                            'Δ'
	'&Dfr;':                             '𝔇'
	'&#120071;':                         '𝔇'
	'&DiacriticalAcute;':                '´'
	'&#180;':                            '´'
	'&DiacriticalDot;':                  '˙'
	'&#729;':                            '˙'
	'&DiacriticalDoubleAcute;':          '˝'
	'&#733;':                            '˝'
	'&DiacriticalGrave;':                '`'
	'&#96;':                             '`'
	'&DiacriticalTilde;':                '˜'
	'&#732;':                            '˜'
	'&Diamond;':                         '⋄'
	'&#8900;':                           '⋄'
	'&DifferentialD;':                   'ⅆ'
	'&#8518;':                           'ⅆ'
	'&Dopf;':                            '𝔻'
	'&#120123;':                         '𝔻'
	'&Dot;':                             '¨'
	'&#168;':                            '¨'
	'&DotDot;':                          '⃜'
	'&#8412;':                           '⃜'
	'&DotEqual;':                        '≐'
	'&#8784;':                           '≐'
	'&DoubleContourIntegral;':           '∯'
	'&DoubleDot;':                       '¨'
	'&DoubleDownArrow;':                 '⇓'
	'&#8659;':                           '⇓'
	'&DoubleLeftArrow;':                 '⇐'
	'&#8656;':                           '⇐'
	'&DoubleLeftRightArrow;':            '⇔'
	'&#8660;':                           '⇔'
	'&DoubleLeftTee;':                   '⫤'
	'&DoubleLongLeftArrow;':             '⟸'
	'&#10232;':                          '⟸'
	'&DoubleLongLeftRightArrow;':        '⟺'
	'&#10234;':                          '⟺'
	'&DoubleLongRightArrow;':            '⟹'
	'&#10233;':                          '⟹'
	'&DoubleRightArrow;':                '⇒'
	'&#8658;':                           '⇒'
	'&DoubleRightTee;':                  '⊨'
	'&#8872;':                           '⊨'
	'&DoubleUpArrow;':                   '⇑'
	'&#8657;':                           '⇑'
	'&DoubleUpDownArrow;':               '⇕'
	'&#8661;':                           '⇕'
	'&DoubleVerticalBar;':               '∥'
	'&#8741;':                           '∥'
	'&DownArrow;':                       '↓'
	'&#8595;':                           '↓'
	'&DownArrowBar;':                    '⤓'
	'&#10515;':                          '⤓'
	'&DownArrowUpArrow;':                '⇵'
	'&#8693;':                           '⇵'
	'&DownBreve;':                       '̑'
	'&#785;':                            '̑'
	'&DownLeftRightVector;':             '⥐'
	'&#10576;':                          '⥐'
	'&DownLeftTeeVector;':               '⥞'
	'&#10590;':                          '⥞'
	'&DownLeftVector;':                  '↽'
	'&#8637;':                           '↽'
	'&DownLeftVectorBar;':               '⥖'
	'&#10582;':                          '⥖'
	'&DownRightTeeVector;':              '⥟'
	'&#10591;':                          '⥟'
	'&DownRightVector;':                 '⇁'
	'&#8641;':                           '⇁'
	'&DownRightVectorBar;':              '⥗'
	'&#10583;':                          '⥗'
	'&DownTee;':                         '⊤'
	'&#8868;':                           '⊤'
	'&DownTeeArrow;':                    '↧'
	'&#8615;':                           '↧'
	'&Downarrow;':                       '⇓'
	'&Dscr;':                            '𝒟'
	'&#119967;':                         '𝒟'
	'&Dstrok;':                          'Đ'
	'&#272;':                            'Đ'
	'&ENG;':                             'Ŋ'
	'&#330;':                            'Ŋ'
	'&#208;':                            'Ð'
	'&ETH;':                             'Ð'
	'&#201;':                            'É'
	'&Eacute;':                          'É'
	'&Ecaron;':                          'Ě'
	'&#282;':                            'Ě'
	'&#202;':                            'Ê'
	'&Ecirc;':                           'Ê'
	'&Ecy;':                             'Э'
	'&#1069;':                           'Э'
	'&Edot;':                            'Ė'
	'&#278;':                            'Ė'
	'&Efr;':                             '𝔈'
	'&#120072;':                         '𝔈'
	'&#200;':                            'È'
	'&Egrave;':                          'È'
	'&Element;':                         '∈'
	'&#8712;':                           '∈'
	'&Emacr;':                           'Ē'
	'&#274;':                            'Ē'
	'&EmptySmallSquare;':                '◻'
	'&#9723;':                           '◻'
	'&EmptyVerySmallSquare;':            '▫'
	'&#9643;':                           '▫'
	'&Eogon;':                           'Ę'
	'&#280;':                            'Ę'
	'&Eopf;':                            '𝔼'
	'&#120124;':                         '𝔼'
	'&Epsilon;':                         'Ε'
	'&#917;':                            'Ε'
	'&Equal;':                           '⩵'
	'&#10869;':                          '⩵'
	'&EqualTilde;':                      '≂'
	'&#8770;':                           '≂'
	'&Equilibrium;':                     '⇌'
	'&#8652;':                           '⇌'
	'&Escr;':                            'ℰ'
	'&#8496;':                           'ℰ'
	'&Esim;':                            '⩳'
	'&#10867;':                          '⩳'
	'&Eta;':                             'Η'
	'&#919;':                            'Η'
	'&#203;':                            'Ë'
	'&Euml;':                            'Ë'
	'&Exists;':                          '∃'
	'&#8707;':                           '∃'
	'&ExponentialE;':                    'ⅇ'
	'&#8519;':                           'ⅇ'
	'&Fcy;':                             'Ф'
	'&#1060;':                           'Ф'
	'&Ffr;':                             '𝔉'
	'&#120073;':                         '𝔉'
	'&FilledSmallSquare;':               '◼'
	'&#9724;':                           '◼'
	'&FilledVerySmallSquare;':           '▪'
	'&#9642;':                           '▪'
	'&Fopf;':                            '𝔽'
	'&#120125;':                         '𝔽'
	'&ForAll;':                          '∀'
	'&#8704;':                           '∀'
	'&Fouriertrf;':                      'ℱ'
	'&#8497;':                           'ℱ'
	'&Fscr;':                            'ℱ'
	'&GJcy;':                            'Ѓ'
	'&#1027;':                           'Ѓ'
	'&#62;':                             '>'
	'&GT;':                              '>'
	'&Gamma;':                           'Γ'
	'&#915;':                            'Γ'
	'&Gammad;':                          'Ϝ'
	'&#988;':                            'Ϝ'
	'&Gbreve;':                          'Ğ'
	'&#286;':                            'Ğ'
	'&Gcedil;':                          'Ģ'
	'&#290;':                            'Ģ'
	'&Gcirc;':                           'Ĝ'
	'&#284;':                            'Ĝ'
	'&Gcy;':                             'Г'
	'&#1043;':                           'Г'
	'&Gdot;':                            'Ġ'
	'&#288;':                            'Ġ'
	'&Gfr;':                             '𝔊'
	'&#120074;':                         '𝔊'
	'&Gg;':                              '⋙'
	'&#8921;':                           '⋙'
	'&Gopf;':                            '𝔾'
	'&#120126;':                         '𝔾'
	'&GreaterEqual;':                    '≥'
	'&#8805;':                           '≥'
	'&GreaterEqualLess;':                '⋛'
	'&#8923;':                           '⋛'
	'&GreaterFullEqual;':                '≧'
	'&#8807;':                           '≧'
	'&GreaterGreater;':                  '⪢'
	'&#10914;':                          '⪢'
	'&GreaterLess;':                     '≷'
	'&#8823;':                           '≷'
	'&GreaterSlantEqual;':               '⩾'
	'&#10878;':                          '⩾'
	'&GreaterTilde;':                    '≳'
	'&#8819;':                           '≳'
	'&Gscr;':                            '𝒢'
	'&#119970;':                         '𝒢'
	'&Gt;':                              '≫'
	'&#8811;':                           '≫'
	'&HARDcy;':                          'Ъ'
	'&#1066;':                           'Ъ'
	'&Hacek;':                           'ˇ'
	'&#711;':                            'ˇ'
	'&Hat;':                             '^'
	'&#94;':                             '^'
	'&Hcirc;':                           'Ĥ'
	'&#292;':                            'Ĥ'
	'&Hfr;':                             'ℌ'
	'&#8460;':                           'ℌ'
	'&HilbertSpace;':                    'ℋ'
	'&#8459;':                           'ℋ'
	'&Hopf;':                            'ℍ'
	'&#8461;':                           'ℍ'
	'&HorizontalLine;':                  '─'
	'&#9472;':                           '─'
	'&Hscr;':                            'ℋ'
	'&Hstrok;':                          'Ħ'
	'&#294;':                            'Ħ'
	'&HumpDownHump;':                    '≎'
	'&HumpEqual;':                       '≏'
	'&#8783;':                           '≏'
	'&IEcy;':                            'Е'
	'&#1045;':                           'Е'
	'&IJlig;':                           'Ĳ'
	'&#306;':                            'Ĳ'
	'&IOcy;':                            'Ё'
	'&#1025;':                           'Ё'
	'&#205;':                            'Í'
	'&Iacute;':                          'Í'
	'&#206;':                            'Î'
	'&Icirc;':                           'Î'
	'&Icy;':                             'И'
	'&#1048;':                           'И'
	'&Idot;':                            'İ'
	'&#304;':                            'İ'
	'&Ifr;':                             'ℑ'
	'&#8465;':                           'ℑ'
	'&#204;':                            'Ì'
	'&Igrave;':                          'Ì'
	'&Im;':                              'ℑ'
	'&Imacr;':                           'Ī'
	'&#298;':                            'Ī'
	'&ImaginaryI;':                      'ⅈ'
	'&#8520;':                           'ⅈ'
	'&Implies;':                         '⇒'
	'&Int;':                             '∬'
	'&#8748;':                           '∬'
	'&Integral;':                        '∫'
	'&#8747;':                           '∫'
	'&Intersection;':                    '⋂'
	'&#8898;':                           '⋂'
	'&InvisibleComma;':                  '⁣'
	'&#8291;':                           '⁣'
	'&InvisibleTimes;':                  '⁢'
	'&#8290;':                           '⁢'
	'&Iogon;':                           'Į'
	'&#302;':                            'Į'
	'&Iopf;':                            '𝕀'
	'&#120128;':                         '𝕀'
	'&Iota;':                            'Ι'
	'&#921;':                            'Ι'
	'&Iscr;':                            'ℐ'
	'&#8464;':                           'ℐ'
	'&Itilde;':                          'Ĩ'
	'&#296;':                            'Ĩ'
	'&Iukcy;':                           'І'
	'&#1030;':                           'І'
	'&#207;':                            'Ï'
	'&Iuml;':                            'Ï'
	'&Jcirc;':                           'Ĵ'
	'&#308;':                            'Ĵ'
	'&Jcy;':                             'Й'
	'&#1049;':                           'Й'
	'&Jfr;':                             '𝔍'
	'&#120077;':                         '𝔍'
	'&Jopf;':                            '𝕁'
	'&#120129;':                         '𝕁'
	'&Jscr;':                            '𝒥'
	'&#119973;':                         '𝒥'
	'&Jsercy;':                          'Ј'
	'&#1032;':                           'Ј'
	'&Jukcy;':                           'Є'
	'&#1028;':                           'Є'
	'&KHcy;':                            'Х'
	'&#1061;':                           'Х'
	'&KJcy;':                            'Ќ'
	'&#1036;':                           'Ќ'
	'&Kappa;':                           'Κ'
	'&#922;':                            'Κ'
	'&Kcedil;':                          'Ķ'
	'&#310;':                            'Ķ'
	'&Kcy;':                             'К'
	'&#1050;':                           'К'
	'&Kfr;':                             '𝔎'
	'&#120078;':                         '𝔎'
	'&Kopf;':                            '𝕂'
	'&#120130;':                         '𝕂'
	'&Kscr;':                            '𝒦'
	'&#119974;':                         '𝒦'
	'&LJcy;':                            'Љ'
	'&#1033;':                           'Љ'
	'&#60;':                             '<'
	'&LT;':                              '<'
	'&Lacute;':                          'Ĺ'
	'&#313;':                            'Ĺ'
	'&Lambda;':                          'Λ'
	'&#923;':                            'Λ'
	'&Lang;':                            '⟪'
	'&#10218;':                          '⟪'
	'&Laplacetrf;':                      'ℒ'
	'&#8466;':                           'ℒ'
	'&Larr;':                            '↞'
	'&#8606;':                           '↞'
	'&Lcaron;':                          'Ľ'
	'&#317;':                            'Ľ'
	'&Lcedil;':                          'Ļ'
	'&#315;':                            'Ļ'
	'&Lcy;':                             'Л'
	'&#1051;':                           'Л'
	'&LeftAngleBracket;':                '⟨'
	'&#10216;':                          '⟨'
	'&LeftArrow;':                       '←'
	'&#8592;':                           '←'
	'&LeftArrowBar;':                    '⇤'
	'&#8676;':                           '⇤'
	'&LeftArrowRightArrow;':             '⇆'
	'&#8646;':                           '⇆'
	'&LeftCeiling;':                     '⌈'
	'&#8968;':                           '⌈'
	'&LeftDoubleBracket;':               '⟦'
	'&#10214;':                          '⟦'
	'&LeftDownTeeVector;':               '⥡'
	'&#10593;':                          '⥡'
	'&LeftDownVector;':                  '⇃'
	'&#8643;':                           '⇃'
	'&LeftDownVectorBar;':               '⥙'
	'&#10585;':                          '⥙'
	'&LeftFloor;':                       '⌊'
	'&#8970;':                           '⌊'
	'&LeftRightArrow;':                  '↔'
	'&#8596;':                           '↔'
	'&LeftRightVector;':                 '⥎'
	'&#10574;':                          '⥎'
	'&LeftTee;':                         '⊣'
	'&#8867;':                           '⊣'
	'&LeftTeeArrow;':                    '↤'
	'&#8612;':                           '↤'
	'&LeftTeeVector;':                   '⥚'
	'&#10586;':                          '⥚'
	'&LeftTriangle;':                    '⊲'
	'&#8882;':                           '⊲'
	'&LeftTriangleBar;':                 '⧏'
	'&#10703;':                          '⧏'
	'&LeftTriangleEqual;':               '⊴'
	'&#8884;':                           '⊴'
	'&LeftUpDownVector;':                '⥑'
	'&#10577;':                          '⥑'
	'&LeftUpTeeVector;':                 '⥠'
	'&#10592;':                          '⥠'
	'&LeftUpVector;':                    '↿'
	'&#8639;':                           '↿'
	'&LeftUpVectorBar;':                 '⥘'
	'&#10584;':                          '⥘'
	'&LeftVector;':                      '↼'
	'&#8636;':                           '↼'
	'&LeftVectorBar;':                   '⥒'
	'&#10578;':                          '⥒'
	'&Leftarrow;':                       '⇐'
	'&Leftrightarrow;':                  '⇔'
	'&LessEqualGreater;':                '⋚'
	'&#8922;':                           '⋚'
	'&LessFullEqual;':                   '≦'
	'&#8806;':                           '≦'
	'&LessGreater;':                     '≶'
	'&#8822;':                           '≶'
	'&LessLess;':                        '⪡'
	'&#10913;':                          '⪡'
	'&LessSlantEqual;':                  '⩽'
	'&#10877;':                          '⩽'
	'&LessTilde;':                       '≲'
	'&#8818;':                           '≲'
	'&Lfr;':                             '𝔏'
	'&#120079;':                         '𝔏'
	'&Ll;':                              '⋘'
	'&#8920;':                           '⋘'
	'&Lleftarrow;':                      '⇚'
	'&#8666;':                           '⇚'
	'&Lmidot;':                          'Ŀ'
	'&#319;':                            'Ŀ'
	'&LongLeftArrow;':                   '⟵'
	'&#10229;':                          '⟵'
	'&LongLeftRightArrow;':              '⟷'
	'&#10231;':                          '⟷'
	'&LongRightArrow;':                  '⟶'
	'&#10230;':                          '⟶'
	'&Longleftarrow;':                   '⟸'
	'&Longleftrightarrow;':              '⟺'
	'&Longrightarrow;':                  '⟹'
	'&Lopf;':                            '𝕃'
	'&#120131;':                         '𝕃'
	'&LowerLeftArrow;':                  '↙'
	'&#8601;':                           '↙'
	'&LowerRightArrow;':                 '↘'
	'&#8600;':                           '↘'
	'&Lscr;':                            'ℒ'
	'&Lsh;':                             '↰'
	'&#8624;':                           '↰'
	'&Lstrok;':                          'Ł'
	'&#321;':                            'Ł'
	'&Lt;':                              '≪'
	'&#8810;':                           '≪'
	'&Map;':                             '⤅'
	'&#10501;':                          '⤅'
	'&Mcy;':                             'М'
	'&#1052;':                           'М'
	'&MediumSpace;':                     ' '
	'&#8287;':                           ' '
	'&Mellintrf;':                       'ℳ'
	'&#8499;':                           'ℳ'
	'&Mfr;':                             '𝔐'
	'&#120080;':                         '𝔐'
	'&MinusPlus;':                       '∓'
	'&#8723;':                           '∓'
	'&Mopf;':                            '𝕄'
	'&#120132;':                         '𝕄'
	'&Mscr;':                            'ℳ'
	'&Mu;':                              'Μ'
	'&#924;':                            'Μ'
	'&NJcy;':                            'Њ'
	'&#1034;':                           'Њ'
	'&Nacute;':                          'Ń'
	'&#323;':                            'Ń'
	'&Ncaron;':                          'Ň'
	'&#327;':                            'Ň'
	'&Ncedil;':                          'Ņ'
	'&#325;':                            'Ņ'
	'&Ncy;':                             'Н'
	'&#1053;':                           'Н'
	'&NegativeMediumSpace;':             '​'
	'&#8203;':                           '​'
	'&NegativeThickSpace;':              '​'
	'&NegativeThinSpace;':               '​'
	'&NegativeVeryThinSpace;':           '​'
	'&NestedGreaterGreater;':            '≫'
	'&NestedLessLess;':                  '≪'
	'&NewLine;':                         ''
	'&#10;':                             ''
	'&Nfr;':                             '𝔑'
	'&#120081;':                         '𝔑'
	'&NoBreak;':                         '⁠'
	'&#8288;':                           '⁠'
	'&NonBreakingSpace;':                ' '
	'&#160;':                            ' '
	'&Nopf;':                            'ℕ'
	'&#8469;':                           'ℕ'
	'&Not;':                             '⫬'
	'&#10988;':                          '⫬'
	'&NotCongruent;':                    '≢'
	'&#8802;':                           '≢'
	'&NotCupCap;':                       '≭'
	'&#8813;':                           '≭'
	'&NotDoubleVerticalBar;':            '∦'
	'&#8742;':                           '∦'
	'&NotElement;':                      '∉'
	'&#8713;':                           '∉'
	'&NotEqual;':                        '≠'
	'&#8800;':                           '≠'
	'&NotEqualTilde;':                   '≂'
	'&#8770, 824;':                      '≂'
	'&NotExists;':                       '∄'
	'&#8708;':                           '∄'
	'&NotGreater;':                      '≯'
	'&#8815;':                           '≯'
	'&NotGreaterEqual;':                 '≱'
	'&#8817;':                           '≱'
	'&NotGreaterFullEqual;':             '≧'
	'&#8807, 824;':                      '≧'
	'&NotGreaterGreater;':               '≫'
	'&#8811, 824;':                      '≫'
	'&NotGreaterLess;':                  '≹'
	'&#8825;':                           '≹'
	'&NotGreaterSlantEqual;':            '⩾'
	'&#10878, 824;':                     '⩾'
	'&NotGreaterTilde;':                 '≵'
	'&#8821;':                           '≵'
	'&NotHumpDownHump;':                 '≎'
	'&#8782, 824;':                      '≎'
	'&NotHumpEqual;':                    '≏'
	'&#8783, 824;':                      '≏'
	'&NotLeftTriangle;':                 '⋪'
	'&#8938;':                           '⋪'
	'&NotLeftTriangleBar;':              '⧏'
	'&#10703, 824;':                     '⧏'
	'&NotLeftTriangleEqual;':            '⋬'
	'&#8940;':                           '⋬'
	'&NotLess;':                         '≮'
	'&#8814;':                           '≮'
	'&NotLessEqual;':                    '≰'
	'&#8816;':                           '≰'
	'&NotLessGreater;':                  '≸'
	'&#8824;':                           '≸'
	'&NotLessLess;':                     '≪'
	'&#8810, 824;':                      '≪'
	'&NotLessSlantEqual;':               '⩽'
	'&#10877, 824;':                     '⩽'
	'&NotLessTilde;':                    '≴'
	'&#8820;':                           '≴'
	'&NotNestedGreaterGreater;':         '⪢'
	'&#10914, 824;':                     '⪢'
	'&NotNestedLessLess;':               '⪡'
	'&#10913, 824;':                     '⪡'
	'&NotPrecedes;':                     '⊀'
	'&#8832;':                           '⊀'
	'&NotPrecedesEqual;':                '⪯'
	'&#10927, 824;':                     '⪯'
	'&NotPrecedesSlantEqual;':           '⋠'
	'&#8928;':                           '⋠'
	'&NotReverseElement;':               '∌'
	'&#8716;':                           '∌'
	'&NotRightTriangle;':                '⋫'
	'&#8939;':                           '⋫'
	'&NotRightTriangleBar;':             '⧐'
	'&#10704, 824;':                     '⧐'
	'&NotRightTriangleEqual;':           '⋭'
	'&#8941;':                           '⋭'
	'&NotSquareSubset;':                 '⊏'
	'&#8847, 824;':                      '⊏'
	'&NotSquareSubsetEqual;':            '⋢'
	'&#8930;':                           '⋢'
	'&NotSquareSuperset;':               '⊐'
	'&#8848, 824;':                      '⊐'
	'&NotSquareSupersetEqual;':          '⋣'
	'&#8931;':                           '⋣'
	'&NotSubset;':                       '⊂'
	'&#8834, 8402;':                     '⊂'
	'&NotSubsetEqual;':                  '⊈'
	'&#8840;':                           '⊈'
	'&NotSucceeds;':                     '⊁'
	'&#8833;':                           '⊁'
	'&NotSucceedsEqual;':                '⪰'
	'&#10928, 824;':                     '⪰'
	'&NotSucceedsSlantEqual;':           '⋡'
	'&#8929;':                           '⋡'
	'&NotSucceedsTilde;':                '≿'
	'&#8831, 824;':                      '≿'
	'&NotSuperset;':                     '⊃'
	'&#8835, 8402;':                     '⊃'
	'&NotSupersetEqual;':                '⊉'
	'&#8841;':                           '⊉'
	'&NotTilde;':                        '≁'
	'&#8769;':                           '≁'
	'&NotTildeEqual;':                   '≄'
	'&#8772;':                           '≄'
	'&NotTildeFullEqual;':               '≇'
	'&#8775;':                           '≇'
	'&NotTildeTilde;':                   '≉'
	'&#8777;':                           '≉'
	'&NotVerticalBar;':                  '∤'
	'&#8740;':                           '∤'
	'&Nscr;':                            '𝒩'
	'&#119977;':                         '𝒩'
	'&#209;':                            'Ñ'
	'&Ntilde;':                          'Ñ'
	'&Nu;':                              'Ν'
	'&#925;':                            'Ν'
	'&OElig;':                           'Œ'
	'&#338;':                            'Œ'
	'&#211;':                            'Ó'
	'&Oacute;':                          'Ó'
	'&#212;':                            'Ô'
	'&Ocirc;':                           'Ô'
	'&Ocy;':                             'О'
	'&#1054;':                           'О'
	'&Odblac;':                          'Ő'
	'&#336;':                            'Ő'
	'&Ofr;':                             '𝔒'
	'&#120082;':                         '𝔒'
	'&#210;':                            'Ò'
	'&Ograve;':                          'Ò'
	'&Omacr;':                           'Ō'
	'&#332;':                            'Ō'
	'&Omega;':                           'Ω'
	'&#937;':                            'Ω'
	'&Omicron;':                         'Ο'
	'&#927;':                            'Ο'
	'&Oopf;':                            '𝕆'
	'&#120134;':                         '𝕆'
	'&OpenCurlyDoubleQuote;':            '“'
	'&#8220;':                           '“'
	'&OpenCurlyQuote;':                  '‘'
	'&#8216;':                           '‘'
	'&Or;':                              '⩔'
	'&#10836;':                          '⩔'
	'&Oscr;':                            '𝒪'
	'&#119978;':                         '𝒪'
	'&#216;':                            'Ø'
	'&Oslash;':                          'Ø'
	'&#213;':                            'Õ'
	'&Otilde;':                          'Õ'
	'&Otimes;':                          '⨷'
	'&#10807;':                          '⨷'
	'&#214;':                            'Ö'
	'&Ouml;':                            'Ö'
	'&OverBar;':                         '‾'
	'&#8254;':                           '‾'
	'&OverBrace;':                       '⏞'
	'&#9182;':                           '⏞'
	'&OverBracket;':                     '⎴'
	'&#9140;':                           '⎴'
	'&OverParenthesis;':                 '⏜'
	'&#9180;':                           '⏜'
	'&PartialD;':                        '∂'
	'&#8706;':                           '∂'
	'&Pcy;':                             'П'
	'&#1055;':                           'П'
	'&Pfr;':                             '𝔓'
	'&#120083;':                         '𝔓'
	'&Phi;':                             'Φ'
	'&#934;':                            'Φ'
	'&Pi;':                              'Π'
	'&#928;':                            'Π'
	'&PlusMinus;':                       '±'
	'&#177;':                            '±'
	'&Poincareplane;':                   'ℌ'
	'&Popf;':                            'ℙ'
	'&#8473;':                           'ℙ'
	'&Pr;':                              '⪻'
	'&#10939;':                          '⪻'
	'&Precedes;':                        '≺'
	'&#8826;':                           '≺'
	'&PrecedesEqual;':                   '⪯'
	'&#10927;':                          '⪯'
	'&PrecedesSlantEqual;':              '≼'
	'&#8828;':                           '≼'
	'&PrecedesTilde;':                   '≾'
	'&#8830;':                           '≾'
	'&Prime;':                           '″'
	'&#8243;':                           '″'
	'&Product;':                         '∏'
	'&#8719;':                           '∏'
	'&Proportion;':                      '∷'
	'&Proportional;':                    '∝'
	'&#8733;':                           '∝'
	'&Pscr;':                            '𝒫'
	'&#119979;':                         '𝒫'
	'&Psi;':                             'Ψ'
	'&#936;':                            'Ψ'
	'&#34;':                             '"'
	'&QUOT;':                            '"'
	'&Qfr;':                             '𝔔'
	'&#120084;':                         '𝔔'
	'&Qopf;':                            'ℚ'
	'&#8474;':                           'ℚ'
	'&Qscr;':                            '𝒬'
	'&#119980;':                         '𝒬'
	'&RBarr;':                           '⤐'
	'&#10512;':                          '⤐'
	'&#174;':                            '®'
	'&REG;':                             '®'
	'&Racute;':                          'Ŕ'
	'&#340;':                            'Ŕ'
	'&Rang;':                            '⟫'
	'&#10219;':                          '⟫'
	'&Rarr;':                            '↠'
	'&#8608;':                           '↠'
	'&Rarrtl;':                          '⤖'
	'&#10518;':                          '⤖'
	'&Rcaron;':                          'Ř'
	'&#344;':                            'Ř'
	'&Rcedil;':                          'Ŗ'
	'&#342;':                            'Ŗ'
	'&Rcy;':                             'Р'
	'&#1056;':                           'Р'
	'&Re;':                              'ℜ'
	'&#8476;':                           'ℜ'
	'&ReverseElement;':                  '∋'
	'&#8715;':                           '∋'
	'&ReverseEquilibrium;':              '⇋'
	'&#8651;':                           '⇋'
	'&ReverseUpEquilibrium;':            '⥯'
	'&#10607;':                          '⥯'
	'&Rfr;':                             'ℜ'
	'&Rho;':                             'Ρ'
	'&#929;':                            'Ρ'
	'&RightAngleBracket;':               '⟩'
	'&#10217;':                          '⟩'
	'&RightArrow;':                      '→'
	'&#8594;':                           '→'
	'&RightArrowBar;':                   '⇥'
	'&#8677;':                           '⇥'
	'&RightArrowLeftArrow;':             '⇄'
	'&#8644;':                           '⇄'
	'&RightCeiling;':                    '⌉'
	'&#8969;':                           '⌉'
	'&RightDoubleBracket;':              '⟧'
	'&#10215;':                          '⟧'
	'&RightDownTeeVector;':              '⥝'
	'&#10589;':                          '⥝'
	'&RightDownVector;':                 '⇂'
	'&#8642;':                           '⇂'
	'&RightDownVectorBar;':              '⥕'
	'&#10581;':                          '⥕'
	'&RightFloor;':                      '⌋'
	'&#8971;':                           '⌋'
	'&RightTee;':                        '⊢'
	'&#8866;':                           '⊢'
	'&RightTeeArrow;':                   '↦'
	'&#8614;':                           '↦'
	'&RightTeeVector;':                  '⥛'
	'&#10587;':                          '⥛'
	'&RightTriangle;':                   '⊳'
	'&#8883;':                           '⊳'
	'&RightTriangleBar;':                '⧐'
	'&#10704;':                          '⧐'
	'&RightTriangleEqual;':              '⊵'
	'&#8885;':                           '⊵'
	'&RightUpDownVector;':               '⥏'
	'&#10575;':                          '⥏'
	'&RightUpTeeVector;':                '⥜'
	'&#10588;':                          '⥜'
	'&RightUpVector;':                   '↾'
	'&#8638;':                           '↾'
	'&RightUpVectorBar;':                '⥔'
	'&#10580;':                          '⥔'
	'&RightVector;':                     '⇀'
	'&#8640;':                           '⇀'
	'&RightVectorBar;':                  '⥓'
	'&#10579;':                          '⥓'
	'&Rightarrow;':                      '⇒'
	'&Ropf;':                            'ℝ'
	'&#8477;':                           'ℝ'
	'&RoundImplies;':                    '⥰'
	'&#10608;':                          '⥰'
	'&Rrightarrow;':                     '⇛'
	'&#8667;':                           '⇛'
	'&Rscr;':                            'ℛ'
	'&#8475;':                           'ℛ'
	'&Rsh;':                             '↱'
	'&#8625;':                           '↱'
	'&RuleDelayed;':                     '⧴'
	'&#10740;':                          '⧴'
	'&SHCHcy;':                          'Щ'
	'&#1065;':                           'Щ'
	'&SHcy;':                            'Ш'
	'&#1064;':                           'Ш'
	'&SOFTcy;':                          'Ь'
	'&#1068;':                           'Ь'
	'&Sacute;':                          'Ś'
	'&#346;':                            'Ś'
	'&Sc;':                              '⪼'
	'&#10940;':                          '⪼'
	'&Scaron;':                          'Š'
	'&#352;':                            'Š'
	'&Scedil;':                          'Ş'
	'&#350;':                            'Ş'
	'&Scirc;':                           'Ŝ'
	'&#348;':                            'Ŝ'
	'&Scy;':                             'С'
	'&#1057;':                           'С'
	'&Sfr;':                             '𝔖'
	'&#120086;':                         '𝔖'
	'&ShortDownArrow;':                  '↓'
	'&ShortLeftArrow;':                  '←'
	'&ShortRightArrow;':                 '→'
	'&ShortUpArrow;':                    '↑'
	'&#8593;':                           '↑'
	'&Sigma;':                           'Σ'
	'&#931;':                            'Σ'
	'&SmallCircle;':                     '∘'
	'&#8728;':                           '∘'
	'&Sopf;':                            '𝕊'
	'&#120138;':                         '𝕊'
	'&Sqrt;':                            '√'
	'&#8730;':                           '√'
	'&Square;':                          '□'
	'&#9633;':                           '□'
	'&SquareIntersection;':              '⊓'
	'&#8851;':                           '⊓'
	'&SquareSubset;':                    '⊏'
	'&#8847;':                           '⊏'
	'&SquareSubsetEqual;':               '⊑'
	'&#8849;':                           '⊑'
	'&SquareSuperset;':                  '⊐'
	'&#8848;':                           '⊐'
	'&SquareSupersetEqual;':             '⊒'
	'&#8850;':                           '⊒'
	'&SquareUnion;':                     '⊔'
	'&#8852;':                           '⊔'
	'&Sscr;':                            '𝒮'
	'&#119982;':                         '𝒮'
	'&Star;':                            '⋆'
	'&#8902;':                           '⋆'
	'&Sub;':                             '⋐'
	'&#8912;':                           '⋐'
	'&Subset;':                          '⋐'
	'&SubsetEqual;':                     '⊆'
	'&#8838;':                           '⊆'
	'&Succeeds;':                        '≻'
	'&#8827;':                           '≻'
	'&SucceedsEqual;':                   '⪰'
	'&#10928;':                          '⪰'
	'&SucceedsSlantEqual;':              '≽'
	'&#8829;':                           '≽'
	'&SucceedsTilde;':                   '≿'
	'&#8831;':                           '≿'
	'&SuchThat;':                        '∋'
	'&Sum;':                             '∑'
	'&#8721;':                           '∑'
	'&Sup;':                             '⋑'
	'&#8913;':                           '⋑'
	'&Superset;':                        '⊃'
	'&#8835;':                           '⊃'
	'&SupersetEqual;':                   '⊇'
	'&#8839;':                           '⊇'
	'&Supset;':                          '⋑'
	'&#222;':                            'Þ'
	'&THORN;':                           'Þ'
	'&TRADE;':                           '™'
	'&#8482;':                           '™'
	'&TSHcy;':                           'Ћ'
	'&#1035;':                           'Ћ'
	'&TScy;':                            'Ц'
	'&#1062;':                           'Ц'
	'&Tab;':                             '	'
	'&#9;':                              '	'
	'&Tau;':                             'Τ'
	'&#932;':                            'Τ'
	'&Tcaron;':                          'Ť'
	'&#356;':                            'Ť'
	'&Tcedil;':                          'Ţ'
	'&#354;':                            'Ţ'
	'&Tcy;':                             'Т'
	'&#1058;':                           'Т'
	'&Tfr;':                             '𝔗'
	'&#120087;':                         '𝔗'
	'&Therefore;':                       '∴'
	'&#8756;':                           '∴'
	'&Theta;':                           'Θ'
	'&#920;':                            'Θ'
	'&ThickSpace;':                      ' '
	'&#8287, 8202;':                     ' '
	'&ThinSpace;':                       ' '
	'&#8201;':                           ' '
	'&Tilde;':                           '∼'
	'&#8764;':                           '∼'
	'&TildeEqual;':                      '≃'
	'&#8771;':                           '≃'
	'&TildeFullEqual;':                  '≅'
	'&#8773;':                           '≅'
	'&TildeTilde;':                      '≈'
	'&#8776;':                           '≈'
	'&Topf;':                            '𝕋'
	'&#120139;':                         '𝕋'
	'&TripleDot;':                       '⃛'
	'&#8411;':                           '⃛'
	'&Tscr;':                            '𝒯'
	'&#119983;':                         '𝒯'
	'&Tstrok;':                          'Ŧ'
	'&#358;':                            'Ŧ'
	'&#218;':                            'Ú'
	'&Uacute;':                          'Ú'
	'&Uarr;':                            '↟'
	'&#8607;':                           '↟'
	'&Uarrocir;':                        '⥉'
	'&#10569;':                          '⥉'
	'&Ubrcy;':                           'Ў'
	'&#1038;':                           'Ў'
	'&Ubreve;':                          'Ŭ'
	'&#364;':                            'Ŭ'
	'&#219;':                            'Û'
	'&Ucirc;':                           'Û'
	'&Ucy;':                             'У'
	'&#1059;':                           'У'
	'&Udblac;':                          'Ű'
	'&#368;':                            'Ű'
	'&Ufr;':                             '𝔘'
	'&#120088;':                         '𝔘'
	'&#217;':                            'Ù'
	'&Ugrave;':                          'Ù'
	'&Umacr;':                           'Ū'
	'&#362;':                            'Ū'
	'&UnderBar;':                        '_'
	'&#95;':                             '_'
	'&UnderBrace;':                      '⏟'
	'&#9183;':                           '⏟'
	'&UnderBracket;':                    '⎵'
	'&#9141;':                           '⎵'
	'&UnderParenthesis;':                '⏝'
	'&#9181;':                           '⏝'
	'&Union;':                           '⋃'
	'&#8899;':                           '⋃'
	'&UnionPlus;':                       '⊎'
	'&#8846;':                           '⊎'
	'&Uogon;':                           'Ų'
	'&#370;':                            'Ų'
	'&Uopf;':                            '𝕌'
	'&#120140;':                         '𝕌'
	'&UpArrow;':                         '↑'
	'&UpArrowBar;':                      '⤒'
	'&#10514;':                          '⤒'
	'&UpArrowDownArrow;':                '⇅'
	'&#8645;':                           '⇅'
	'&UpDownArrow;':                     '↕'
	'&#8597;':                           '↕'
	'&UpEquilibrium;':                   '⥮'
	'&#10606;':                          '⥮'
	'&UpTee;':                           '⊥'
	'&#8869;':                           '⊥'
	'&UpTeeArrow;':                      '↥'
	'&#8613;':                           '↥'
	'&Uparrow;':                         '⇑'
	'&Updownarrow;':                     '⇕'
	'&UpperLeftArrow;':                  '↖'
	'&#8598;':                           '↖'
	'&UpperRightArrow;':                 '↗'
	'&#8599;':                           '↗'
	'&Upsi;':                            'ϒ'
	'&#978;':                            'ϒ'
	'&Upsilon;':                         'Υ'
	'&#933;':                            'Υ'
	'&Uring;':                           'Ů'
	'&#366;':                            'Ů'
	'&Uscr;':                            '𝒰'
	'&#119984;':                         '𝒰'
	'&Utilde;':                          'Ũ'
	'&#360;':                            'Ũ'
	'&#220;':                            'Ü'
	'&Uuml;':                            'Ü'
	'&VDash;':                           '⊫'
	'&#8875;':                           '⊫'
	'&Vbar;':                            '⫫'
	'&#10987;':                          '⫫'
	'&Vcy;':                             'В'
	'&#1042;':                           'В'
	'&Vdash;':                           '⊩'
	'&#8873;':                           '⊩'
	'&Vdashl;':                          '⫦'
	'&#10982;':                          '⫦'
	'&Vee;':                             '⋁'
	'&#8897;':                           '⋁'
	'&Verbar;':                          '‖'
	'&#8214;':                           '‖'
	'&Vert;':                            '‖'
	'&VerticalBar;':                     '∣'
	'&#8739;':                           '∣'
	'&VerticalLine;':                    '|'
	'&#124;':                            '|'
	'&VerticalSeparator;':               '❘'
	'&#10072;':                          '❘'
	'&VerticalTilde;':                   '≀'
	'&#8768;':                           '≀'
	'&VeryThinSpace;':                   ' '
	'&#8202;':                           ' '
	'&Vfr;':                             '𝔙'
	'&#120089;':                         '𝔙'
	'&Vopf;':                            '𝕍'
	'&#120141;':                         '𝕍'
	'&Vscr;':                            '𝒱'
	'&#119985;':                         '𝒱'
	'&Vvdash;':                          '⊪'
	'&#8874;':                           '⊪'
	'&Wcirc;':                           'Ŵ'
	'&#372;':                            'Ŵ'
	'&Wedge;':                           '⋀'
	'&#8896;':                           '⋀'
	'&Wfr;':                             '𝔚'
	'&#120090;':                         '𝔚'
	'&Wopf;':                            '𝕎'
	'&#120142;':                         '𝕎'
	'&Wscr;':                            '𝒲'
	'&#119986;':                         '𝒲'
	'&Xfr;':                             '𝔛'
	'&#120091;':                         '𝔛'
	'&Xi;':                              'Ξ'
	'&#926;':                            'Ξ'
	'&Xopf;':                            '𝕏'
	'&#120143;':                         '𝕏'
	'&Xscr;':                            '𝒳'
	'&#119987;':                         '𝒳'
	'&YAcy;':                            'Я'
	'&#1071;':                           'Я'
	'&YIcy;':                            'Ї'
	'&#1031;':                           'Ї'
	'&YUcy;':                            'Ю'
	'&#1070;':                           'Ю'
	'&#221;':                            'Ý'
	'&Yacute;':                          'Ý'
	'&Ycirc;':                           'Ŷ'
	'&#374;':                            'Ŷ'
	'&Ycy;':                             'Ы'
	'&#1067;':                           'Ы'
	'&Yfr;':                             '𝔜'
	'&#120092;':                         '𝔜'
	'&Yopf;':                            '𝕐'
	'&#120144;':                         '𝕐'
	'&Yscr;':                            '𝒴'
	'&#119988;':                         '𝒴'
	'&Yuml;':                            'Ÿ'
	'&#376;':                            'Ÿ'
	'&ZHcy;':                            'Ж'
	'&#1046;':                           'Ж'
	'&Zacute;':                          'Ź'
	'&#377;':                            'Ź'
	'&Zcaron;':                          'Ž'
	'&#381;':                            'Ž'
	'&Zcy;':                             'З'
	'&#1047;':                           'З'
	'&Zdot;':                            'Ż'
	'&#379;':                            'Ż'
	'&ZeroWidthSpace;':                  '​'
	'&Zeta;':                            'Ζ'
	'&#918;':                            'Ζ'
	'&Zfr;':                             'ℨ'
	'&#8488;':                           'ℨ'
	'&Zopf;':                            'ℤ'
	'&#8484;':                           'ℤ'
	'&Zscr;':                            '𝒵'
	'&#119989;':                         '𝒵'
	'&#225;':                            'á'
	'&aacute;':                          'á'
	'&abreve;':                          'ă'
	'&#259;':                            'ă'
	'&ac;':                              '∾'
	'&#8766;':                           '∾'
	'&acE;':                             '∾'
	'&#8766, 819;':                      '∾'
	'&acd;':                             '∿'
	'&#8767;':                           '∿'
	'&#226;':                            'â'
	'&acirc;':                           'â'
	'&acute;':                           '´'
	'&acy;':                             'а'
	'&#1072;':                           'а'
	'&#230;':                            'æ'
	'&aelig;':                           'æ'
	'&af;':                              '⁡'
	'&afr;':                             '𝔞'
	'&#120094;':                         '𝔞'
	'&#224;':                            'à'
	'&agrave;':                          'à'
	'&alefsym;':                         'ℵ'
	'&#8501;':                           'ℵ'
	'&aleph;':                           'ℵ'
	'&alpha;':                           'α'
	'&#945;':                            'α'
	'&amacr;':                           'ā'
	'&#257;':                            'ā'
	'&amalg;':                           '⨿'
	'&#10815;':                          '⨿'
	'&amp;':                             '&'
	'&and;':                             '∧'
	'&#8743;':                           '∧'
	'&andand;':                          '⩕'
	'&#10837;':                          '⩕'
	'&andd;':                            '⩜'
	'&#10844;':                          '⩜'
	'&andslope;':                        '⩘'
	'&#10840;':                          '⩘'
	'&andv;':                            '⩚'
	'&#10842;':                          '⩚'
	'&ang;':                             '∠'
	'&#8736;':                           '∠'
	'&ange;':                            '⦤'
	'&#10660;':                          '⦤'
	'&angle;':                           '∠'
	'&angmsd;':                          '∡'
	'&#8737;':                           '∡'
	'&angmsdaa;':                        '⦨'
	'&#10664;':                          '⦨'
	'&angmsdab;':                        '⦩'
	'&#10665;':                          '⦩'
	'&angmsdac;':                        '⦪'
	'&#10666;':                          '⦪'
	'&angmsdad;':                        '⦫'
	'&#10667;':                          '⦫'
	'&angmsdae;':                        '⦬'
	'&#10668;':                          '⦬'
	'&angmsdaf;':                        '⦭'
	'&#10669;':                          '⦭'
	'&angmsdag;':                        '⦮'
	'&#10670;':                          '⦮'
	'&angmsdah;':                        '⦯'
	'&#10671;':                          '⦯'
	'&angrt;':                           '∟'
	'&#8735;':                           '∟'
	'&angrtvb;':                         '⊾'
	'&#8894;':                           '⊾'
	'&angrtvbd;':                        '⦝'
	'&#10653;':                          '⦝'
	'&angsph;':                          '∢'
	'&#8738;':                           '∢'
	'&angst;':                           'Å'
	'&angzarr;':                         '⍼'
	'&#9084;':                           '⍼'
	'&aogon;':                           'ą'
	'&#261;':                            'ą'
	'&aopf;':                            '𝕒'
	'&#120146;':                         '𝕒'
	'&ap;':                              '≈'
	'&apE;':                             '⩰'
	'&#10864;':                          '⩰'
	'&apacir;':                          '⩯'
	'&#10863;':                          '⩯'
	'&ape;':                             '≊'
	'&#8778;':                           '≊'
	'&apid;':                            '≋'
	'&#8779;':                           '≋'
	'&apos;':                            "'"
	'&#39;':                             "'"
	'&approx;':                          '≈'
	'&approxeq;':                        '≊'
	'&#229;':                            'å'
	'&aring;':                           'å'
	'&ascr;':                            '𝒶'
	'&#119990;':                         '𝒶'
	'&ast;':                             '*'
	'&#42;':                             '*'
	'&asymp;':                           '≈'
	'&asympeq;':                         '≍'
	'&#227;':                            'ã'
	'&atilde;':                          'ã'
	'&#228;':                            'ä'
	'&auml;':                            'ä'
	'&awconint;':                        '∳'
	'&awint;':                           '⨑'
	'&#10769;':                          '⨑'
	'&bNot;':                            '⫭'
	'&#10989;':                          '⫭'
	'&backcong;':                        '≌'
	'&#8780;':                           '≌'
	'&backepsilon;':                     '϶'
	'&#1014;':                           '϶'
	'&backprime;':                       '‵'
	'&#8245;':                           '‵'
	'&backsim;':                         '∽'
	'&#8765;':                           '∽'
	'&backsimeq;':                       '⋍'
	'&#8909;':                           '⋍'
	'&barvee;':                          '⊽'
	'&#8893;':                           '⊽'
	'&barwed;':                          '⌅'
	'&#8965;':                           '⌅'
	'&barwedge;':                        '⌅'
	'&bbrk;':                            '⎵'
	'&bbrktbrk;':                        '⎶'
	'&#9142;':                           '⎶'
	'&bcong;':                           '≌'
	'&bcy;':                             'б'
	'&#1073;':                           'б'
	'&bdquo;':                           '„'
	'&#8222;':                           '„'
	'&becaus;':                          '∵'
	'&because;':                         '∵'
	'&bemptyv;':                         '⦰'
	'&#10672;':                          '⦰'
	'&bepsi;':                           '϶'
	'&bernou;':                          'ℬ'
	'&beta;':                            'β'
	'&#946;':                            'β'
	'&beth;':                            'ℶ'
	'&#8502;':                           'ℶ'
	'&between;':                         '≬'
	'&#8812;':                           '≬'
	'&bfr;':                             '𝔟'
	'&#120095;':                         '𝔟'
	'&bigcap;':                          '⋂'
	'&bigcirc;':                         '◯'
	'&#9711;':                           '◯'
	'&bigcup;':                          '⋃'
	'&bigodot;':                         '⨀'
	'&#10752;':                          '⨀'
	'&bigoplus;':                        '⨁'
	'&#10753;':                          '⨁'
	'&bigotimes;':                       '⨂'
	'&#10754;':                          '⨂'
	'&bigsqcup;':                        '⨆'
	'&#10758;':                          '⨆'
	'&bigstar;':                         '★'
	'&#9733;':                           '★'
	'&bigtriangledown;':                 '▽'
	'&#9661;':                           '▽'
	'&bigtriangleup;':                   '△'
	'&#9651;':                           '△'
	'&biguplus;':                        '⨄'
	'&#10756;':                          '⨄'
	'&bigvee;':                          '⋁'
	'&bigwedge;':                        '⋀'
	'&bkarow;':                          '⤍'
	'&#10509;':                          '⤍'
	'&blacklozenge;':                    '⧫'
	'&#10731;':                          '⧫'
	'&blacksquare;':                     '▪'
	'&blacktriangle;':                   '▴'
	'&#9652;':                           '▴'
	'&blacktriangledown;':               '▾'
	'&#9662;':                           '▾'
	'&blacktriangleleft;':               '◂'
	'&#9666;':                           '◂'
	'&blacktriangleright;':              '▸'
	'&#9656;':                           '▸'
	'&blank;':                           '␣'
	'&#9251;':                           '␣'
	'&blk12;':                           '▒'
	'&#9618;':                           '▒'
	'&blk14;':                           '░'
	'&#9617;':                           '░'
	'&blk34;':                           '▓'
	'&#9619;':                           '▓'
	'&block;':                           '█'
	'&#9608;':                           '█'
	'&bne;':                             '='
	'&#61, 8421;':                       '='
	'&bnequiv;':                         '≡'
	'&#8801, 8421;':                     '≡'
	'&bnot;':                            '⌐'
	'&#8976;':                           '⌐'
	'&bopf;':                            '𝕓'
	'&#120147;':                         '𝕓'
	'&bot;':                             '⊥'
	'&bottom;':                          '⊥'
	'&bowtie;':                          '⋈'
	'&#8904;':                           '⋈'
	'&boxDL;':                           '╗'
	'&#9559;':                           '╗'
	'&boxDR;':                           '╔'
	'&#9556;':                           '╔'
	'&boxDl;':                           '╖'
	'&#9558;':                           '╖'
	'&boxDr;':                           '╓'
	'&#9555;':                           '╓'
	'&boxH;':                            '═'
	'&#9552;':                           '═'
	'&boxHD;':                           '╦'
	'&#9574;':                           '╦'
	'&boxHU;':                           '╩'
	'&#9577;':                           '╩'
	'&boxHd;':                           '╤'
	'&#9572;':                           '╤'
	'&boxHu;':                           '╧'
	'&#9575;':                           '╧'
	'&boxUL;':                           '╝'
	'&#9565;':                           '╝'
	'&boxUR;':                           '╚'
	'&#9562;':                           '╚'
	'&boxUl;':                           '╜'
	'&#9564;':                           '╜'
	'&boxUr;':                           '╙'
	'&#9561;':                           '╙'
	'&boxV;':                            '║'
	'&#9553;':                           '║'
	'&boxVH;':                           '╬'
	'&#9580;':                           '╬'
	'&boxVL;':                           '╣'
	'&#9571;':                           '╣'
	'&boxVR;':                           '╠'
	'&#9568;':                           '╠'
	'&boxVh;':                           '╫'
	'&#9579;':                           '╫'
	'&boxVl;':                           '╢'
	'&#9570;':                           '╢'
	'&boxVr;':                           '╟'
	'&#9567;':                           '╟'
	'&boxbox;':                          '⧉'
	'&#10697;':                          '⧉'
	'&boxdL;':                           '╕'
	'&#9557;':                           '╕'
	'&boxdR;':                           '╒'
	'&#9554;':                           '╒'
	'&boxdl;':                           '┐'
	'&#9488;':                           '┐'
	'&boxdr;':                           '┌'
	'&#9484;':                           '┌'
	'&boxh;':                            '─'
	'&boxhD;':                           '╥'
	'&#9573;':                           '╥'
	'&boxhU;':                           '╨'
	'&#9576;':                           '╨'
	'&boxhd;':                           '┬'
	'&#9516;':                           '┬'
	'&boxhu;':                           '┴'
	'&#9524;':                           '┴'
	'&boxminus;':                        '⊟'
	'&#8863;':                           '⊟'
	'&boxplus;':                         '⊞'
	'&#8862;':                           '⊞'
	'&boxtimes;':                        '⊠'
	'&#8864;':                           '⊠'
	'&boxuL;':                           '╛'
	'&#9563;':                           '╛'
	'&boxuR;':                           '╘'
	'&#9560;':                           '╘'
	'&boxul;':                           '┘'
	'&#9496;':                           '┘'
	'&boxur;':                           '└'
	'&#9492;':                           '└'
	'&boxv;':                            '│'
	'&#9474;':                           '│'
	'&boxvH;':                           '╪'
	'&#9578;':                           '╪'
	'&boxvL;':                           '╡'
	'&#9569;':                           '╡'
	'&boxvR;':                           '╞'
	'&#9566;':                           '╞'
	'&boxvh;':                           '┼'
	'&#9532;':                           '┼'
	'&boxvl;':                           '┤'
	'&#9508;':                           '┤'
	'&boxvr;':                           '├'
	'&#9500;':                           '├'
	'&bprime;':                          '‵'
	'&breve;':                           '˘'
	'&#166;':                            '¦'
	'&brvbar;':                          '¦'
	'&bscr;':                            '𝒷'
	'&#119991;':                         '𝒷'
	'&bsemi;':                           '⁏'
	'&#8271;':                           '⁏'
	'&bsim;':                            '∽'
	'&bsime;':                           '⋍'
	'&bsol;':                            '\\'
	'&#92;':                             '\\'
	'&bsolb;':                           '⧅'
	'&#10693;':                          '⧅'
	'&bsolhsub;':                        '⟈'
	'&#10184;':                          '⟈'
	'&bull;':                            '•'
	'&#8226;':                           '•'
	'&bullet;':                          '•'
	'&bump;':                            '≎'
	'&bumpE;':                           '⪮'
	'&#10926;':                          '⪮'
	'&bumpe;':                           '≏'
	'&bumpeq;':                          '≏'
	'&cacute;':                          'ć'
	'&#263;':                            'ć'
	'&cap;':                             '∩'
	'&#8745;':                           '∩'
	'&capand;':                          '⩄'
	'&#10820;':                          '⩄'
	'&capbrcup;':                        '⩉'
	'&#10825;':                          '⩉'
	'&capcap;':                          '⩋'
	'&#10827;':                          '⩋'
	'&capcup;':                          '⩇'
	'&#10823;':                          '⩇'
	'&capdot;':                          '⩀'
	'&#10816;':                          '⩀'
	'&caps;':                            '∩'
	'&#8745, 65024;':                    '∩'
	'&caret;':                           '⁁'
	'&#8257;':                           '⁁'
	'&caron;':                           'ˇ'
	'&ccaps;':                           '⩍'
	'&#10829;':                          '⩍'
	'&ccaron;':                          'č'
	'&#269;':                            'č'
	'&#231;':                            'ç'
	'&ccedil;':                          'ç'
	'&ccirc;':                           'ĉ'
	'&#265;':                            'ĉ'
	'&ccups;':                           '⩌'
	'&#10828;':                          '⩌'
	'&ccupssm;':                         '⩐'
	'&#10832;':                          '⩐'
	'&cdot;':                            'ċ'
	'&#267;':                            'ċ'
	'&cedil;':                           '¸'
	'&cemptyv;':                         '⦲'
	'&#10674;':                          '⦲'
	'&#162;':                            '¢'
	'&cent;':                            '¢'
	'&centerdot;':                       '·'
	'&cfr;':                             '𝔠'
	'&#120096;':                         '𝔠'
	'&chcy;':                            'ч'
	'&#1095;':                           'ч'
	'&check;':                           '✓'
	'&#10003;':                          '✓'
	'&checkmark;':                       '✓'
	'&chi;':                             'χ'
	'&#967;':                            'χ'
	'&cir;':                             '○'
	'&#9675;':                           '○'
	'&cirE;':                            '⧃'
	'&#10691;':                          '⧃'
	'&circ;':                            'ˆ'
	'&#710;':                            'ˆ'
	'&circeq;':                          '≗'
	'&#8791;':                           '≗'
	'&circlearrowleft;':                 '↺'
	'&#8634;':                           '↺'
	'&circlearrowright;':                '↻'
	'&#8635;':                           '↻'
	'&circledR;':                        '®'
	'&circledS;':                        'Ⓢ'
	'&#9416;':                           'Ⓢ'
	'&circledast;':                      '⊛'
	'&#8859;':                           '⊛'
	'&circledcirc;':                     '⊚'
	'&#8858;':                           '⊚'
	'&circleddash;':                     '⊝'
	'&#8861;':                           '⊝'
	'&cire;':                            '≗'
	'&cirfnint;':                        '⨐'
	'&#10768;':                          '⨐'
	'&cirmid;':                          '⫯'
	'&#10991;':                          '⫯'
	'&cirscir;':                         '⧂'
	'&#10690;':                          '⧂'
	'&clubs;':                           '♣'
	'&#9827;':                           '♣'
	'&clubsuit;':                        '♣'
	'&colon;':                           ':'
	'&#58;':                             ':'
	'&colone;':                          '≔'
	'&coloneq;':                         '≔'
	'&comma;':                           ','
	'&#44;':                             ','
	'&commat;':                          '@'
	'&#64;':                             '@'
	'&comp;':                            '∁'
	'&#8705;':                           '∁'
	'&compfn;':                          '∘'
	'&complement;':                      '∁'
	'&complexes;':                       'ℂ'
	'&cong;':                            '≅'
	'&congdot;':                         '⩭'
	'&#10861;':                          '⩭'
	'&conint;':                          '∮'
	'&copf;':                            '𝕔'
	'&#120148;':                         '𝕔'
	'&coprod;':                          '∐'
	'&copy;':                            '©'
	'&copysr;':                          '℗'
	'&#8471;':                           '℗'
	'&crarr;':                           '↵'
	'&#8629;':                           '↵'
	'&cross;':                           '✗'
	'&#10007;':                          '✗'
	'&cscr;':                            '𝒸'
	'&#119992;':                         '𝒸'
	'&csub;':                            '⫏'
	'&#10959;':                          '⫏'
	'&csube;':                           '⫑'
	'&#10961;':                          '⫑'
	'&csup;':                            '⫐'
	'&#10960;':                          '⫐'
	'&csupe;':                           '⫒'
	'&#10962;':                          '⫒'
	'&ctdot;':                           '⋯'
	'&#8943;':                           '⋯'
	'&cudarrl;':                         '⤸'
	'&#10552;':                          '⤸'
	'&cudarrr;':                         '⤵'
	'&#10549;':                          '⤵'
	'&cuepr;':                           '⋞'
	'&#8926;':                           '⋞'
	'&cuesc;':                           '⋟'
	'&#8927;':                           '⋟'
	'&cularr;':                          '↶'
	'&#8630;':                           '↶'
	'&cularrp;':                         '⤽'
	'&#10557;':                          '⤽'
	'&cup;':                             '∪'
	'&#8746;':                           '∪'
	'&cupbrcap;':                        '⩈'
	'&#10824;':                          '⩈'
	'&cupcap;':                          '⩆'
	'&#10822;':                          '⩆'
	'&cupcup;':                          '⩊'
	'&#10826;':                          '⩊'
	'&cupdot;':                          '⊍'
	'&#8845;':                           '⊍'
	'&cupor;':                           '⩅'
	'&#10821;':                          '⩅'
	'&cups;':                            '∪'
	'&#8746, 65024;':                    '∪'
	'&curarr;':                          '↷'
	'&#8631;':                           '↷'
	'&curarrm;':                         '⤼'
	'&#10556;':                          '⤼'
	'&curlyeqprec;':                     '⋞'
	'&curlyeqsucc;':                     '⋟'
	'&curlyvee;':                        '⋎'
	'&#8910;':                           '⋎'
	'&curlywedge;':                      '⋏'
	'&#8911;':                           '⋏'
	'&#164;':                            '¤'
	'&curren;':                          '¤'
	'&curvearrowleft;':                  '↶'
	'&curvearrowright;':                 '↷'
	'&cuvee;':                           '⋎'
	'&cuwed;':                           '⋏'
	'&cwconint;':                        '∲'
	'&cwint;':                           '∱'
	'&#8753;':                           '∱'
	'&cylcty;':                          '⌭'
	'&#9005;':                           '⌭'
	'&dArr;':                            '⇓'
	'&dHar;':                            '⥥'
	'&#10597;':                          '⥥'
	'&dagger;':                          '†'
	'&#8224;':                           '†'
	'&daleth;':                          'ℸ'
	'&#8504;':                           'ℸ'
	'&darr;':                            '↓'
	'&dash;':                            '‐'
	'&#8208;':                           '‐'
	'&dashv;':                           '⊣'
	'&dbkarow;':                         '⤏'
	'&#10511;':                          '⤏'
	'&dblac;':                           '˝'
	'&dcaron;':                          'ď'
	'&#271;':                            'ď'
	'&dcy;':                             'д'
	'&#1076;':                           'д'
	'&dd;':                              'ⅆ'
	'&ddagger;':                         '‡'
	'&ddarr;':                           '⇊'
	'&#8650;':                           '⇊'
	'&ddotseq;':                         '⩷'
	'&#10871;':                          '⩷'
	'&#176;':                            '°'
	'&deg;':                             '°'
	'&delta;':                           'δ'
	'&#948;':                            'δ'
	'&demptyv;':                         '⦱'
	'&#10673;':                          '⦱'
	'&dfisht;':                          '⥿'
	'&#10623;':                          '⥿'
	'&dfr;':                             '𝔡'
	'&#120097;':                         '𝔡'
	'&dharl;':                           '⇃'
	'&dharr;':                           '⇂'
	'&diam;':                            '⋄'
	'&diamond;':                         '⋄'
	'&diamondsuit;':                     '♦'
	'&#9830;':                           '♦'
	'&diams;':                           '♦'
	'&die;':                             '¨'
	'&digamma;':                         'ϝ'
	'&#989;':                            'ϝ'
	'&disin;':                           '⋲'
	'&#8946;':                           '⋲'
	'&div;':                             '÷'
	'&#247;':                            '÷'
	'&divide;':                          '÷'
	'&divideontimes;':                   '⋇'
	'&#8903;':                           '⋇'
	'&divonx;':                          '⋇'
	'&djcy;':                            'ђ'
	'&#1106;':                           'ђ'
	'&dlcorn;':                          '⌞'
	'&#8990;':                           '⌞'
	'&dlcrop;':                          '⌍'
	'&#8973;':                           '⌍'
	'&dollar;':                          '$'
	'&#36;':                             '$'
	'&dopf;':                            '𝕕'
	'&#120149;':                         '𝕕'
	'&dot;':                             '˙'
	'&doteq;':                           '≐'
	'&doteqdot;':                        '≑'
	'&#8785;':                           '≑'
	'&dotminus;':                        '∸'
	'&#8760;':                           '∸'
	'&dotplus;':                         '∔'
	'&#8724;':                           '∔'
	'&dotsquare;':                       '⊡'
	'&#8865;':                           '⊡'
	'&doublebarwedge;':                  '⌆'
	'&downarrow;':                       '↓'
	'&downdownarrows;':                  '⇊'
	'&downharpoonleft;':                 '⇃'
	'&downharpoonright;':                '⇂'
	'&drbkarow;':                        '⤐'
	'&drcorn;':                          '⌟'
	'&#8991;':                           '⌟'
	'&drcrop;':                          '⌌'
	'&#8972;':                           '⌌'
	'&dscr;':                            '𝒹'
	'&#119993;':                         '𝒹'
	'&dscy;':                            'ѕ'
	'&#1109;':                           'ѕ'
	'&dsol;':                            '⧶'
	'&#10742;':                          '⧶'
	'&dstrok;':                          'đ'
	'&#273;':                            'đ'
	'&dtdot;':                           '⋱'
	'&#8945;':                           '⋱'
	'&dtri;':                            '▿'
	'&#9663;':                           '▿'
	'&dtrif;':                           '▾'
	'&duarr;':                           '⇵'
	'&duhar;':                           '⥯'
	'&dwangle;':                         '⦦'
	'&#10662;':                          '⦦'
	'&dzcy;':                            'џ'
	'&#1119;':                           'џ'
	'&dzigrarr;':                        '⟿'
	'&#10239;':                          '⟿'
	'&eDDot;':                           '⩷'
	'&eDot;':                            '≑'
	'&#233;':                            'é'
	'&eacute;':                          'é'
	'&easter;':                          '⩮'
	'&#10862;':                          '⩮'
	'&ecaron;':                          'ě'
	'&#283;':                            'ě'
	'&ecir;':                            '≖'
	'&#8790;':                           '≖'
	'&#234;':                            'ê'
	'&ecirc;':                           'ê'
	'&ecolon;':                          '≕'
	'&#8789;':                           '≕'
	'&ecy;':                             'э'
	'&#1101;':                           'э'
	'&edot;':                            'ė'
	'&#279;':                            'ė'
	'&ee;':                              'ⅇ'
	'&efDot;':                           '≒'
	'&#8786;':                           '≒'
	'&efr;':                             '𝔢'
	'&#120098;':                         '𝔢'
	'&eg;':                              '⪚'
	'&#10906;':                          '⪚'
	'&#232;':                            'è'
	'&egrave;':                          'è'
	'&egs;':                             '⪖'
	'&#10902;':                          '⪖'
	'&egsdot;':                          '⪘'
	'&#10904;':                          '⪘'
	'&el;':                              '⪙'
	'&#10905;':                          '⪙'
	'&elinters;':                        '⏧'
	'&#9191;':                           '⏧'
	'&ell;':                             'ℓ'
	'&#8467;':                           'ℓ'
	'&els;':                             '⪕'
	'&#10901;':                          '⪕'
	'&elsdot;':                          '⪗'
	'&#10903;':                          '⪗'
	'&emacr;':                           'ē'
	'&#275;':                            'ē'
	'&empty;':                           '∅'
	'&#8709;':                           '∅'
	'&emptyset;':                        '∅'
	'&emptyv;':                          '∅'
	'&emsp13;':                          ' '
	'&#8196;':                           ' '
	'&emsp14;':                          ' '
	'&#8197;':                           ' '
	'&emsp;':                            ' '
	'&#8195;':                           ' '
	'&eng;':                             'ŋ'
	'&#331;':                            'ŋ'
	'&ensp;':                            ' '
	'&#8194;':                           ' '
	'&eogon;':                           'ę'
	'&#281;':                            'ę'
	'&eopf;':                            '𝕖'
	'&#120150;':                         '𝕖'
	'&epar;':                            '⋕'
	'&#8917;':                           '⋕'
	'&eparsl;':                          '⧣'
	'&#10723;':                          '⧣'
	'&eplus;':                           '⩱'
	'&#10865;':                          '⩱'
	'&epsi;':                            'ε'
	'&#949;':                            'ε'
	'&epsilon;':                         'ε'
	'&epsiv;':                           'ϵ'
	'&#1013;':                           'ϵ'
	'&eqcirc;':                          '≖'
	'&eqcolon;':                         '≕'
	'&eqsim;':                           '≂'
	'&eqslantgtr;':                      '⪖'
	'&eqslantless;':                     '⪕'
	'&equals;':                          '='
	'&#61;':                             '='
	'&equest;':                          '≟'
	'&#8799;':                           '≟'
	'&equiv;':                           '≡'
	'&equivDD;':                         '⩸'
	'&#10872;':                          '⩸'
	'&eqvparsl;':                        '⧥'
	'&#10725;':                          '⧥'
	'&erDot;':                           '≓'
	'&#8787;':                           '≓'
	'&erarr;':                           '⥱'
	'&#10609;':                          '⥱'
	'&escr;':                            'ℯ'
	'&#8495;':                           'ℯ'
	'&esdot;':                           '≐'
	'&esim;':                            '≂'
	'&eta;':                             'η'
	'&#951;':                            'η'
	'&#240;':                            'ð'
	'&eth;':                             'ð'
	'&#235;':                            'ë'
	'&euml;':                            'ë'
	'&euro;':                            '€'
	'&#8364;':                           '€'
	'&excl;':                            '!'
	'&#33;':                             '!'
	'&exist;':                           '∃'
	'&expectation;':                     'ℰ'
	'&exponentiale;':                    'ⅇ'
	'&fallingdotseq;':                   '≒'
	'&fcy;':                             'ф'
	'&#1092;':                           'ф'
	'&female;':                          '♀'
	'&#9792;':                           '♀'
	'&ffilig;':                          'ﬃ'
	'&#64259;':                          'ﬃ'
	'&fflig;':                           'ﬀ'
	'&#64256;':                          'ﬀ'
	'&ffllig;':                          'ﬄ'
	'&#64260;':                          'ﬄ'
	'&ffr;':                             '𝔣'
	'&#120099;':                         '𝔣'
	'&filig;':                           'ﬁ'
	'&#64257;':                          'ﬁ'
	'&fjlig;':                           'f'
	'&#102, 106;':                       'f'
	'&flat;':                            '♭'
	'&#9837;':                           '♭'
	'&fllig;':                           'ﬂ'
	'&#64258;':                          'ﬂ'
	'&fltns;':                           '▱'
	'&#9649;':                           '▱'
	'&fnof;':                            'ƒ'
	'&#402;':                            'ƒ'
	'&fopf;':                            '𝕗'
	'&#120151;':                         '𝕗'
	'&forall;':                          '∀'
	'&fork;':                            '⋔'
	'&#8916;':                           '⋔'
	'&forkv;':                           '⫙'
	'&#10969;':                          '⫙'
	'&fpartint;':                        '⨍'
	'&#10765;':                          '⨍'
	'&#189;':                            '½'
	'&frac12;':                          '½'
	'&frac13;':                          '⅓'
	'&#8531;':                           '⅓'
	'&#188;':                            '¼'
	'&frac14;':                          '¼'
	'&frac15;':                          '⅕'
	'&#8533;':                           '⅕'
	'&frac16;':                          '⅙'
	'&#8537;':                           '⅙'
	'&frac18;':                          '⅛'
	'&#8539;':                           '⅛'
	'&frac23;':                          '⅔'
	'&#8532;':                           '⅔'
	'&frac25;':                          '⅖'
	'&#8534;':                           '⅖'
	'&#190;':                            '¾'
	'&frac34;':                          '¾'
	'&frac35;':                          '⅗'
	'&#8535;':                           '⅗'
	'&frac38;':                          '⅜'
	'&#8540;':                           '⅜'
	'&frac45;':                          '⅘'
	'&#8536;':                           '⅘'
	'&frac56;':                          '⅚'
	'&#8538;':                           '⅚'
	'&frac58;':                          '⅝'
	'&#8541;':                           '⅝'
	'&frac78;':                          '⅞'
	'&#8542;':                           '⅞'
	'&frasl;':                           '⁄'
	'&#8260;':                           '⁄'
	'&frown;':                           '⌢'
	'&#8994;':                           '⌢'
	'&fscr;':                            '𝒻'
	'&#119995;':                         '𝒻'
	'&gE;':                              '≧'
	'&gEl;':                             '⪌'
	'&#10892;':                          '⪌'
	'&gacute;':                          'ǵ'
	'&#501;':                            'ǵ'
	'&gamma;':                           'γ'
	'&#947;':                            'γ'
	'&gammad;':                          'ϝ'
	'&gap;':                             '⪆'
	'&#10886;':                          '⪆'
	'&gbreve;':                          'ğ'
	'&#287;':                            'ğ'
	'&gcirc;':                           'ĝ'
	'&#285;':                            'ĝ'
	'&gcy;':                             'г'
	'&#1075;':                           'г'
	'&gdot;':                            'ġ'
	'&#289;':                            'ġ'
	'&ge;':                              '≥'
	'&gel;':                             '⋛'
	'&geq;':                             '≥'
	'&geqq;':                            '≧'
	'&geqslant;':                        '⩾'
	'&ges;':                             '⩾'
	'&gescc;':                           '⪩'
	'&#10921;':                          '⪩'
	'&gesdot;':                          '⪀'
	'&#10880;':                          '⪀'
	'&gesdoto;':                         '⪂'
	'&#10882;':                          '⪂'
	'&gesdotol;':                        '⪄'
	'&#10884;':                          '⪄'
	'&gesl;':                            '⋛'
	'&#8923, 65024;':                    '⋛'
	'&gesles;':                          '⪔'
	'&#10900;':                          '⪔'
	'&gfr;':                             '𝔤'
	'&#120100;':                         '𝔤'
	'&gg;':                              '≫'
	'&ggg;':                             '⋙'
	'&gimel;':                           'ℷ'
	'&#8503;':                           'ℷ'
	'&gjcy;':                            'ѓ'
	'&#1107;':                           'ѓ'
	'&gl;':                              '≷'
	'&glE;':                             '⪒'
	'&#10898;':                          '⪒'
	'&gla;':                             '⪥'
	'&#10917;':                          '⪥'
	'&glj;':                             '⪤'
	'&#10916;':                          '⪤'
	'&gnE;':                             '≩'
	'&#8809;':                           '≩'
	'&gnap;':                            '⪊'
	'&#10890;':                          '⪊'
	'&gnapprox;':                        '⪊'
	'&gne;':                             '⪈'
	'&#10888;':                          '⪈'
	'&gneq;':                            '⪈'
	'&gneqq;':                           '≩'
	'&gnsim;':                           '⋧'
	'&#8935;':                           '⋧'
	'&gopf;':                            '𝕘'
	'&#120152;':                         '𝕘'
	'&grave;':                           '`'
	'&gscr;':                            'ℊ'
	'&#8458;':                           'ℊ'
	'&gsim;':                            '≳'
	'&gsime;':                           '⪎'
	'&#10894;':                          '⪎'
	'&gsiml;':                           '⪐'
	'&#10896;':                          '⪐'
	'&gt;':                              '>'
	'&gtcc;':                            '⪧'
	'&#10919;':                          '⪧'
	'&gtcir;':                           '⩺'
	'&#10874;':                          '⩺'
	'&gtdot;':                           '⋗'
	'&#8919;':                           '⋗'
	'&gtlPar;':                          '⦕'
	'&#10645;':                          '⦕'
	'&gtquest;':                         '⩼'
	'&#10876;':                          '⩼'
	'&gtrapprox;':                       '⪆'
	'&gtrarr;':                          '⥸'
	'&#10616;':                          '⥸'
	'&gtrdot;':                          '⋗'
	'&gtreqless;':                       '⋛'
	'&gtreqqless;':                      '⪌'
	'&gtrless;':                         '≷'
	'&gtrsim;':                          '≳'
	'&gvertneqq;':                       '≩'
	'&#8809, 65024;':                    '≩'
	'&gvnE;':                            '≩'
	'&hArr;':                            '⇔'
	'&hairsp;':                          ' '
	'&half;':                            '½'
	'&hamilt;':                          'ℋ'
	'&hardcy;':                          'ъ'
	'&#1098;':                           'ъ'
	'&harr;':                            '↔'
	'&harrcir;':                         '⥈'
	'&#10568;':                          '⥈'
	'&harrw;':                           '↭'
	'&#8621;':                           '↭'
	'&hbar;':                            'ℏ'
	'&#8463;':                           'ℏ'
	'&hcirc;':                           'ĥ'
	'&#293;':                            'ĥ'
	'&hearts;':                          '♥'
	'&#9829;':                           '♥'
	'&heartsuit;':                       '♥'
	'&hellip;':                          '…'
	'&#8230;':                           '…'
	'&hercon;':                          '⊹'
	'&#8889;':                           '⊹'
	'&hfr;':                             '𝔥'
	'&#120101;':                         '𝔥'
	'&hksearow;':                        '⤥'
	'&#10533;':                          '⤥'
	'&hkswarow;':                        '⤦'
	'&#10534;':                          '⤦'
	'&hoarr;':                           '⇿'
	'&#8703;':                           '⇿'
	'&homtht;':                          '∻'
	'&#8763;':                           '∻'
	'&hookleftarrow;':                   '↩'
	'&#8617;':                           '↩'
	'&hookrightarrow;':                  '↪'
	'&#8618;':                           '↪'
	'&hopf;':                            '𝕙'
	'&#120153;':                         '𝕙'
	'&horbar;':                          '―'
	'&#8213;':                           '―'
	'&hscr;':                            '𝒽'
	'&#119997;':                         '𝒽'
	'&hslash;':                          'ℏ'
	'&hstrok;':                          'ħ'
	'&#295;':                            'ħ'
	'&hybull;':                          '⁃'
	'&#8259;':                           '⁃'
	'&hyphen;':                          '‐'
	'&#237;':                            'í'
	'&iacute;':                          'í'
	'&ic;':                              '⁣'
	'&#238;':                            'î'
	'&icirc;':                           'î'
	'&icy;':                             'и'
	'&#1080;':                           'и'
	'&iecy;':                            'е'
	'&#1077;':                           'е'
	'&#161;':                            '¡'
	'&iexcl;':                           '¡'
	'&iff;':                             '⇔'
	'&ifr;':                             '𝔦'
	'&#120102;':                         '𝔦'
	'&#236;':                            'ì'
	'&igrave;':                          'ì'
	'&ii;':                              'ⅈ'
	'&iiiint;':                          '⨌'
	'&#10764;':                          '⨌'
	'&iiint;':                           '∭'
	'&#8749;':                           '∭'
	'&iinfin;':                          '⧜'
	'&#10716;':                          '⧜'
	'&iiota;':                           '℩'
	'&#8489;':                           '℩'
	'&ijlig;':                           'ĳ'
	'&#307;':                            'ĳ'
	'&imacr;':                           'ī'
	'&#299;':                            'ī'
	'&image;':                           'ℑ'
	'&imagline;':                        'ℐ'
	'&imagpart;':                        'ℑ'
	'&imath;':                           'ı'
	'&#305;':                            'ı'
	'&imof;':                            '⊷'
	'&#8887;':                           '⊷'
	'&imped;':                           'Ƶ'
	'&#437;':                            'Ƶ'
	'&in;':                              '∈'
	'&incare;':                          '℅'
	'&#8453;':                           '℅'
	'&infin;':                           '∞'
	'&#8734;':                           '∞'
	'&infintie;':                        '⧝'
	'&#10717;':                          '⧝'
	'&inodot;':                          'ı'
	'&int;':                             '∫'
	'&intcal;':                          '⊺'
	'&#8890;':                           '⊺'
	'&integers;':                        'ℤ'
	'&intercal;':                        '⊺'
	'&intlarhk;':                        '⨗'
	'&#10775;':                          '⨗'
	'&intprod;':                         '⨼'
	'&#10812;':                          '⨼'
	'&iocy;':                            'ё'
	'&#1105;':                           'ё'
	'&iogon;':                           'į'
	'&#303;':                            'į'
	'&iopf;':                            '𝕚'
	'&#120154;':                         '𝕚'
	'&iota;':                            'ι'
	'&#953;':                            'ι'
	'&iprod;':                           '⨼'
	'&#191;':                            '¿'
	'&iquest;':                          '¿'
	'&iscr;':                            '𝒾'
	'&#119998;':                         '𝒾'
	'&isin;':                            '∈'
	'&isinE;':                           '⋹'
	'&#8953;':                           '⋹'
	'&isindot;':                         '⋵'
	'&#8949;':                           '⋵'
	'&isins;':                           '⋴'
	'&#8948;':                           '⋴'
	'&isinsv;':                          '⋳'
	'&#8947;':                           '⋳'
	'&isinv;':                           '∈'
	'&it;':                              '⁢'
	'&itilde;':                          'ĩ'
	'&#297;':                            'ĩ'
	'&iukcy;':                           'і'
	'&#1110;':                           'і'
	'&#239;':                            'ï'
	'&iuml;':                            'ï'
	'&jcirc;':                           'ĵ'
	'&#309;':                            'ĵ'
	'&jcy;':                             'й'
	'&#1081;':                           'й'
	'&jfr;':                             '𝔧'
	'&#120103;':                         '𝔧'
	'&jmath;':                           'ȷ'
	'&#567;':                            'ȷ'
	'&jopf;':                            '𝕛'
	'&#120155;':                         '𝕛'
	'&jscr;':                            '𝒿'
	'&#119999;':                         '𝒿'
	'&jsercy;':                          'ј'
	'&#1112;':                           'ј'
	'&jukcy;':                           'є'
	'&#1108;':                           'є'
	'&kappa;':                           'κ'
	'&#954;':                            'κ'
	'&kappav;':                          'ϰ'
	'&#1008;':                           'ϰ'
	'&kcedil;':                          'ķ'
	'&#311;':                            'ķ'
	'&kcy;':                             'к'
	'&#1082;':                           'к'
	'&kfr;':                             '𝔨'
	'&#120104;':                         '𝔨'
	'&kgreen;':                          'ĸ'
	'&#312;':                            'ĸ'
	'&khcy;':                            'х'
	'&#1093;':                           'х'
	'&kjcy;':                            'ќ'
	'&#1116;':                           'ќ'
	'&kopf;':                            '𝕜'
	'&#120156;':                         '𝕜'
	'&kscr;':                            '𝓀'
	'&#120000;':                         '𝓀'
	'&lAarr;':                           '⇚'
	'&lArr;':                            '⇐'
	'&lAtail;':                          '⤛'
	'&#10523;':                          '⤛'
	'&lBarr;':                           '⤎'
	'&#10510;':                          '⤎'
	'&lE;':                              '≦'
	'&lEg;':                             '⪋'
	'&#10891;':                          '⪋'
	'&lHar;':                            '⥢'
	'&#10594;':                          '⥢'
	'&lacute;':                          'ĺ'
	'&#314;':                            'ĺ'
	'&laemptyv;':                        '⦴'
	'&#10676;':                          '⦴'
	'&lagran;':                          'ℒ'
	'&lambda;':                          'λ'
	'&#955;':                            'λ'
	'&lang;':                            '⟨'
	'&langd;':                           '⦑'
	'&#10641;':                          '⦑'
	'&langle;':                          '⟨'
	'&lap;':                             '⪅'
	'&#10885;':                          '⪅'
	'&#171;':                            '«'
	'&laquo;':                           '«'
	'&larr;':                            '←'
	'&larrb;':                           '⇤'
	'&larrbfs;':                         '⤟'
	'&#10527;':                          '⤟'
	'&larrfs;':                          '⤝'
	'&#10525;':                          '⤝'
	'&larrhk;':                          '↩'
	'&larrlp;':                          '↫'
	'&#8619;':                           '↫'
	'&larrpl;':                          '⤹'
	'&#10553;':                          '⤹'
	'&larrsim;':                         '⥳'
	'&#10611;':                          '⥳'
	'&larrtl;':                          '↢'
	'&#8610;':                           '↢'
	'&lat;':                             '⪫'
	'&#10923;':                          '⪫'
	'&latail;':                          '⤙'
	'&#10521;':                          '⤙'
	'&late;':                            '⪭'
	'&#10925;':                          '⪭'
	'&lates;':                           '⪭'
	'&#10925, 65024;':                   '⪭'
	'&lbarr;':                           '⤌'
	'&#10508;':                          '⤌'
	'&lbbrk;':                           '❲'
	'&#10098;':                          '❲'
	'&lbrace;':                          '{'
	'&#123;':                            '{'
	'&lbrack;':                          '['
	'&#91;':                             '['
	'&lbrke;':                           '⦋'
	'&#10635;':                          '⦋'
	'&lbrksld;':                         '⦏'
	'&#10639;':                          '⦏'
	'&lbrkslu;':                         '⦍'
	'&#10637;':                          '⦍'
	'&lcaron;':                          'ľ'
	'&#318;':                            'ľ'
	'&lcedil;':                          'ļ'
	'&#316;':                            'ļ'
	'&lceil;':                           '⌈'
	'&lcub;':                            '{'
	'&lcy;':                             'л'
	'&#1083;':                           'л'
	'&ldca;':                            '⤶'
	'&#10550;':                          '⤶'
	'&ldquo;':                           '“'
	'&ldquor;':                          '„'
	'&ldrdhar;':                         '⥧'
	'&#10599;':                          '⥧'
	'&ldrushar;':                        '⥋'
	'&#10571;':                          '⥋'
	'&ldsh;':                            '↲'
	'&#8626;':                           '↲'
	'&le;':                              '≤'
	'&#8804;':                           '≤'
	'&leftarrow;':                       '←'
	'&leftarrowtail;':                   '↢'
	'&leftharpoondown;':                 '↽'
	'&leftharpoonup;':                   '↼'
	'&leftleftarrows;':                  '⇇'
	'&#8647;':                           '⇇'
	'&leftrightarrow;':                  '↔'
	'&leftrightarrows;':                 '⇆'
	'&leftrightharpoons;':               '⇋'
	'&leftrightsquigarrow;':             '↭'
	'&leftthreetimes;':                  '⋋'
	'&#8907;':                           '⋋'
	'&leg;':                             '⋚'
	'&leq;':                             '≤'
	'&leqq;':                            '≦'
	'&leqslant;':                        '⩽'
	'&les;':                             '⩽'
	'&lescc;':                           '⪨'
	'&#10920;':                          '⪨'
	'&lesdot;':                          '⩿'
	'&#10879;':                          '⩿'
	'&lesdoto;':                         '⪁'
	'&#10881;':                          '⪁'
	'&lesdotor;':                        '⪃'
	'&#10883;':                          '⪃'
	'&lesg;':                            '⋚'
	'&#8922, 65024;':                    '⋚'
	'&lesges;':                          '⪓'
	'&#10899;':                          '⪓'
	'&lessapprox;':                      '⪅'
	'&lessdot;':                         '⋖'
	'&#8918;':                           '⋖'
	'&lesseqgtr;':                       '⋚'
	'&lesseqqgtr;':                      '⪋'
	'&lessgtr;':                         '≶'
	'&lesssim;':                         '≲'
	'&lfisht;':                          '⥼'
	'&#10620;':                          '⥼'
	'&lfloor;':                          '⌊'
	'&lfr;':                             '𝔩'
	'&#120105;':                         '𝔩'
	'&lg;':                              '≶'
	'&lgE;':                             '⪑'
	'&#10897;':                          '⪑'
	'&lhard;':                           '↽'
	'&lharu;':                           '↼'
	'&lharul;':                          '⥪'
	'&#10602;':                          '⥪'
	'&lhblk;':                           '▄'
	'&#9604;':                           '▄'
	'&ljcy;':                            'љ'
	'&#1113;':                           'љ'
	'&ll;':                              '≪'
	'&llarr;':                           '⇇'
	'&llcorner;':                        '⌞'
	'&llhard;':                          '⥫'
	'&#10603;':                          '⥫'
	'&lltri;':                           '◺'
	'&#9722;':                           '◺'
	'&lmidot;':                          'ŀ'
	'&#320;':                            'ŀ'
	'&lmoust;':                          '⎰'
	'&#9136;':                           '⎰'
	'&lmoustache;':                      '⎰'
	'&lnE;':                             '≨'
	'&#8808;':                           '≨'
	'&lnap;':                            '⪉'
	'&#10889;':                          '⪉'
	'&lnapprox;':                        '⪉'
	'&lne;':                             '⪇'
	'&#10887;':                          '⪇'
	'&lneq;':                            '⪇'
	'&lneqq;':                           '≨'
	'&lnsim;':                           '⋦'
	'&#8934;':                           '⋦'
	'&loang;':                           '⟬'
	'&#10220;':                          '⟬'
	'&loarr;':                           '⇽'
	'&#8701;':                           '⇽'
	'&lobrk;':                           '⟦'
	'&longleftarrow;':                   '⟵'
	'&longleftrightarrow;':              '⟷'
	'&longmapsto;':                      '⟼'
	'&#10236;':                          '⟼'
	'&longrightarrow;':                  '⟶'
	'&looparrowleft;':                   '↫'
	'&looparrowright;':                  '↬'
	'&#8620;':                           '↬'
	'&lopar;':                           '⦅'
	'&#10629;':                          '⦅'
	'&lopf;':                            '𝕝'
	'&#120157;':                         '𝕝'
	'&loplus;':                          '⨭'
	'&#10797;':                          '⨭'
	'&lotimes;':                         '⨴'
	'&#10804;':                          '⨴'
	'&lowast;':                          '∗'
	'&#8727;':                           '∗'
	'&lowbar;':                          '_'
	'&loz;':                             '◊'
	'&#9674;':                           '◊'
	'&lozenge;':                         '◊'
	'&lozf;':                            '⧫'
	'&lpar;':                            '('
	'&#40;':                             '('
	'&lparlt;':                          '⦓'
	'&#10643;':                          '⦓'
	'&lrarr;':                           '⇆'
	'&lrcorner;':                        '⌟'
	'&lrhar;':                           '⇋'
	'&lrhard;':                          '⥭'
	'&#10605;':                          '⥭'
	'&lrm;':                             '‎'
	'&#8206;':                           '‎'
	'&lrtri;':                           '⊿'
	'&#8895;':                           '⊿'
	'&lsaquo;':                          '‹'
	'&#8249;':                           '‹'
	'&lscr;':                            '𝓁'
	'&#120001;':                         '𝓁'
	'&lsh;':                             '↰'
	'&lsim;':                            '≲'
	'&lsime;':                           '⪍'
	'&#10893;':                          '⪍'
	'&lsimg;':                           '⪏'
	'&#10895;':                          '⪏'
	'&lsqb;':                            '['
	'&lsquo;':                           '‘'
	'&lsquor;':                          '‚'
	'&#8218;':                           '‚'
	'&lstrok;':                          'ł'
	'&#322;':                            'ł'
	'&lt;':                              '<'
	'&ltcc;':                            '⪦'
	'&#10918;':                          '⪦'
	'&ltcir;':                           '⩹'
	'&#10873;':                          '⩹'
	'&ltdot;':                           '⋖'
	'&lthree;':                          '⋋'
	'&ltimes;':                          '⋉'
	'&#8905;':                           '⋉'
	'&ltlarr;':                          '⥶'
	'&#10614;':                          '⥶'
	'&ltquest;':                         '⩻'
	'&#10875;':                          '⩻'
	'&ltrPar;':                          '⦖'
	'&#10646;':                          '⦖'
	'&ltri;':                            '◃'
	'&#9667;':                           '◃'
	'&ltrie;':                           '⊴'
	'&ltrif;':                           '◂'
	'&lurdshar;':                        '⥊'
	'&#10570;':                          '⥊'
	'&luruhar;':                         '⥦'
	'&#10598;':                          '⥦'
	'&lvertneqq;':                       '≨'
	'&#8808, 65024;':                    '≨'
	'&lvnE;':                            '≨'
	'&mDDot;':                           '∺'
	'&#8762;':                           '∺'
	'&#175;':                            '¯'
	'&macr;':                            '¯'
	'&male;':                            '♂'
	'&#9794;':                           '♂'
	'&malt;':                            '✠'
	'&#10016;':                          '✠'
	'&maltese;':                         '✠'
	'&map;':                             '↦'
	'&mapsto;':                          '↦'
	'&mapstodown;':                      '↧'
	'&mapstoleft;':                      '↤'
	'&mapstoup;':                        '↥'
	'&marker;':                          '▮'
	'&#9646;':                           '▮'
	'&mcomma;':                          '⨩'
	'&#10793;':                          '⨩'
	'&mcy;':                             'м'
	'&#1084;':                           'м'
	'&mdash;':                           '—'
	'&#8212;':                           '—'
	'&measuredangle;':                   '∡'
	'&mfr;':                             '𝔪'
	'&#120106;':                         '𝔪'
	'&mho;':                             '℧'
	'&#8487;':                           '℧'
	'&#181;':                            'µ'
	'&micro;':                           'µ'
	'&mid;':                             '∣'
	'&midast;':                          '*'
	'&midcir;':                          '⫰'
	'&#10992;':                          '⫰'
	'&middot;':                          '·'
	'&minus;':                           '−'
	'&#8722;':                           '−'
	'&minusb;':                          '⊟'
	'&minusd;':                          '∸'
	'&minusdu;':                         '⨪'
	'&#10794;':                          '⨪'
	'&mlcp;':                            '⫛'
	'&#10971;':                          '⫛'
	'&mldr;':                            '…'
	'&mnplus;':                          '∓'
	'&models;':                          '⊧'
	'&#8871;':                           '⊧'
	'&mopf;':                            '𝕞'
	'&#120158;':                         '𝕞'
	'&mp;':                              '∓'
	'&mscr;':                            '𝓂'
	'&#120002;':                         '𝓂'
	'&mstpos;':                          '∾'
	'&mu;':                              'μ'
	'&#956;':                            'μ'
	'&multimap;':                        '⊸'
	'&#8888;':                           '⊸'
	'&mumap;':                           '⊸'
	'&nGg;':                             '⋙'
	'&#8921, 824;':                      '⋙'
	'&nGt;':                             '≫'
	'&#8811, 8402;':                     '≫'
	'&nGtv;':                            '≫'
	'&nLeftarrow;':                      '⇍'
	'&#8653;':                           '⇍'
	'&nLeftrightarrow;':                 '⇎'
	'&#8654;':                           '⇎'
	'&nLl;':                             '⋘'
	'&#8920, 824;':                      '⋘'
	'&nLt;':                             '≪'
	'&#8810, 8402;':                     '≪'
	'&nLtv;':                            '≪'
	'&nRightarrow;':                     '⇏'
	'&#8655;':                           '⇏'
	'&nVDash;':                          '⊯'
	'&#8879;':                           '⊯'
	'&nVdash;':                          '⊮'
	'&#8878;':                           '⊮'
	'&nabla;':                           '∇'
	'&nacute;':                          'ń'
	'&#324;':                            'ń'
	'&nang;':                            '∠'
	'&#8736, 8402;':                     '∠'
	'&nap;':                             '≉'
	'&napE;':                            '⩰'
	'&#10864, 824;':                     '⩰'
	'&napid;':                           '≋'
	'&#8779, 824;':                      '≋'
	'&napos;':                           'ŉ'
	'&#329;':                            'ŉ'
	'&napprox;':                         '≉'
	'&natur;':                           '♮'
	'&#9838;':                           '♮'
	'&natural;':                         '♮'
	'&naturals;':                        'ℕ'
	'&nbsp;':                            ' '
	'&nbump;':                           '≎'
	'&nbumpe;':                          '≏'
	'&ncap;':                            '⩃'
	'&#10819;':                          '⩃'
	'&ncaron;':                          'ň'
	'&#328;':                            'ň'
	'&ncedil;':                          'ņ'
	'&#326;':                            'ņ'
	'&ncong;':                           '≇'
	'&ncongdot;':                        '⩭'
	'&#10861, 824;':                     '⩭'
	'&ncup;':                            '⩂'
	'&#10818;':                          '⩂'
	'&ncy;':                             'н'
	'&#1085;':                           'н'
	'&ndash;':                           '–'
	'&#8211;':                           '–'
	'&ne;':                              '≠'
	'&neArr;':                           '⇗'
	'&#8663;':                           '⇗'
	'&nearhk;':                          '⤤'
	'&#10532;':                          '⤤'
	'&nearr;':                           '↗'
	'&nearrow;':                         '↗'
	'&nedot;':                           '≐'
	'&#8784, 824;':                      '≐'
	'&nequiv;':                          '≢'
	'&nesear;':                          '⤨'
	'&#10536;':                          '⤨'
	'&nesim;':                           '≂'
	'&nexist;':                          '∄'
	'&nexists;':                         '∄'
	'&nfr;':                             '𝔫'
	'&#120107;':                         '𝔫'
	'&ngE;':                             '≧'
	'&nge;':                             '≱'
	'&ngeq;':                            '≱'
	'&ngeqq;':                           '≧'
	'&ngeqslant;':                       '⩾'
	'&nges;':                            '⩾'
	'&ngsim;':                           '≵'
	'&ngt;':                             '≯'
	'&ngtr;':                            '≯'
	'&nhArr;':                           '⇎'
	'&nharr;':                           '↮'
	'&#8622;':                           '↮'
	'&nhpar;':                           '⫲'
	'&#10994;':                          '⫲'
	'&ni;':                              '∋'
	'&nis;':                             '⋼'
	'&#8956;':                           '⋼'
	'&nisd;':                            '⋺'
	'&#8954;':                           '⋺'
	'&niv;':                             '∋'
	'&njcy;':                            'њ'
	'&#1114;':                           'њ'
	'&nlArr;':                           '⇍'
	'&nlE;':                             '≦'
	'&#8806, 824;':                      '≦'
	'&nlarr;':                           '↚'
	'&#8602;':                           '↚'
	'&nldr;':                            '‥'
	'&#8229;':                           '‥'
	'&nle;':                             '≰'
	'&nleftarrow;':                      '↚'
	'&nleftrightarrow;':                 '↮'
	'&nleq;':                            '≰'
	'&nleqq;':                           '≦'
	'&nleqslant;':                       '⩽'
	'&nles;':                            '⩽'
	'&nless;':                           '≮'
	'&nlsim;':                           '≴'
	'&nlt;':                             '≮'
	'&nltri;':                           '⋪'
	'&nltrie;':                          '⋬'
	'&nmid;':                            '∤'
	'&nopf;':                            '𝕟'
	'&#120159;':                         '𝕟'
	'&#172;':                            '¬'
	'&not;':                             '¬'
	'&notin;':                           '∉'
	'&notinE;':                          '⋹'
	'&#8953, 824;':                      '⋹'
	'&notindot;':                        '⋵'
	'&#8949, 824;':                      '⋵'
	'&notinva;':                         '∉'
	'&notinvb;':                         '⋷'
	'&#8951;':                           '⋷'
	'&notinvc;':                         '⋶'
	'&#8950;':                           '⋶'
	'&notni;':                           '∌'
	'&notniva;':                         '∌'
	'&notnivb;':                         '⋾'
	'&#8958;':                           '⋾'
	'&notnivc;':                         '⋽'
	'&#8957;':                           '⋽'
	'&npar;':                            '∦'
	'&nparallel;':                       '∦'
	'&nparsl;':                          '⫽'
	'&#11005, 8421;':                    '⫽'
	'&npart;':                           '∂'
	'&#8706, 824;':                      '∂'
	'&npolint;':                         '⨔'
	'&#10772;':                          '⨔'
	'&npr;':                             '⊀'
	'&nprcue;':                          '⋠'
	'&npre;':                            '⪯'
	'&nprec;':                           '⊀'
	'&npreceq;':                         '⪯'
	'&nrArr;':                           '⇏'
	'&nrarr;':                           '↛'
	'&#8603;':                           '↛'
	'&nrarrc;':                          '⤳'
	'&#10547, 824;':                     '⤳'
	'&nrarrw;':                          '↝'
	'&#8605, 824;':                      '↝'
	'&nrightarrow;':                     '↛'
	'&nrtri;':                           '⋫'
	'&nrtrie;':                          '⋭'
	'&nsc;':                             '⊁'
	'&nsccue;':                          '⋡'
	'&nsce;':                            '⪰'
	'&nscr;':                            '𝓃'
	'&#120003;':                         '𝓃'
	'&nshortmid;':                       '∤'
	'&nshortparallel;':                  '∦'
	'&nsim;':                            '≁'
	'&nsime;':                           '≄'
	'&nsimeq;':                          '≄'
	'&nsmid;':                           '∤'
	'&nspar;':                           '∦'
	'&nsqsube;':                         '⋢'
	'&nsqsupe;':                         '⋣'
	'&nsub;':                            '⊄'
	'&#8836;':                           '⊄'
	'&nsubE;':                           '⫅'
	'&#10949, 824;':                     '⫅'
	'&nsube;':                           '⊈'
	'&nsubset;':                         '⊂'
	'&nsubseteq;':                       '⊈'
	'&nsubseteqq;':                      '⫅'
	'&nsucc;':                           '⊁'
	'&nsucceq;':                         '⪰'
	'&nsup;':                            '⊅'
	'&#8837;':                           '⊅'
	'&nsupE;':                           '⫆'
	'&#10950, 824;':                     '⫆'
	'&nsupe;':                           '⊉'
	'&nsupset;':                         '⊃'
	'&nsupseteq;':                       '⊉'
	'&nsupseteqq;':                      '⫆'
	'&ntgl;':                            '≹'
	'&#241;':                            'ñ'
	'&ntilde;':                          'ñ'
	'&ntlg;':                            '≸'
	'&ntriangleleft;':                   '⋪'
	'&ntrianglelefteq;':                 '⋬'
	'&ntriangleright;':                  '⋫'
	'&ntrianglerighteq;':                '⋭'
	'&nu;':                              'ν'
	'&#957;':                            'ν'
	'&num;':                             '#'
	'&#35;':                             '#'
	'&numero;':                          '№'
	'&#8470;':                           '№'
	'&numsp;':                           ' '
	'&#8199;':                           ' '
	'&nvDash;':                          '⊭'
	'&#8877;':                           '⊭'
	'&nvHarr;':                          '⤄'
	'&#10500;':                          '⤄'
	'&nvap;':                            '≍'
	'&#8781, 8402;':                     '≍'
	'&nvdash;':                          '⊬'
	'&#8876;':                           '⊬'
	'&nvge;':                            '≥'
	'&#8805, 8402;':                     '≥'
	'&nvgt;':                            '>'
	'&#62, 8402;':                       '>'
	'&nvinfin;':                         '⧞'
	'&#10718;':                          '⧞'
	'&nvlArr;':                          '⤂'
	'&#10498;':                          '⤂'
	'&nvle;':                            '≤'
	'&#8804, 8402;':                     '≤'
	'&nvlt;':                            '<'
	'&#60, 8402;':                       '<'
	'&nvltrie;':                         '⊴'
	'&#8884, 8402;':                     '⊴'
	'&nvrArr;':                          '⤃'
	'&#10499;':                          '⤃'
	'&nvrtrie;':                         '⊵'
	'&#8885, 8402;':                     '⊵'
	'&nvsim;':                           '∼'
	'&#8764, 8402;':                     '∼'
	'&nwArr;':                           '⇖'
	'&#8662;':                           '⇖'
	'&nwarhk;':                          '⤣'
	'&#10531;':                          '⤣'
	'&nwarr;':                           '↖'
	'&nwarrow;':                         '↖'
	'&nwnear;':                          '⤧'
	'&#10535;':                          '⤧'
	'&oS;':                              'Ⓢ'
	'&#243;':                            'ó'
	'&oacute;':                          'ó'
	'&oast;':                            '⊛'
	'&ocir;':                            '⊚'
	'&#244;':                            'ô'
	'&ocirc;':                           'ô'
	'&ocy;':                             'о'
	'&#1086;':                           'о'
	'&odash;':                           '⊝'
	'&odblac;':                          'ő'
	'&#337;':                            'ő'
	'&odiv;':                            '⨸'
	'&#10808;':                          '⨸'
	'&odot;':                            '⊙'
	'&odsold;':                          '⦼'
	'&#10684;':                          '⦼'
	'&oelig;':                           'œ'
	'&#339;':                            'œ'
	'&ofcir;':                           '⦿'
	'&#10687;':                          '⦿'
	'&ofr;':                             '𝔬'
	'&#120108;':                         '𝔬'
	'&ogon;':                            '˛'
	'&#731;':                            '˛'
	'&#242;':                            'ò'
	'&ograve;':                          'ò'
	'&ogt;':                             '⧁'
	'&#10689;':                          '⧁'
	'&ohbar;':                           '⦵'
	'&#10677;':                          '⦵'
	'&ohm;':                             'Ω'
	'&oint;':                            '∮'
	'&olarr;':                           '↺'
	'&olcir;':                           '⦾'
	'&#10686;':                          '⦾'
	'&olcross;':                         '⦻'
	'&#10683;':                          '⦻'
	'&oline;':                           '‾'
	'&olt;':                             '⧀'
	'&#10688;':                          '⧀'
	'&omacr;':                           'ō'
	'&#333;':                            'ō'
	'&omega;':                           'ω'
	'&#969;':                            'ω'
	'&omicron;':                         'ο'
	'&#959;':                            'ο'
	'&omid;':                            '⦶'
	'&#10678;':                          '⦶'
	'&ominus;':                          '⊖'
	'&oopf;':                            '𝕠'
	'&#120160;':                         '𝕠'
	'&opar;':                            '⦷'
	'&#10679;':                          '⦷'
	'&operp;':                           '⦹'
	'&#10681;':                          '⦹'
	'&oplus;':                           '⊕'
	'&or;':                              '∨'
	'&#8744;':                           '∨'
	'&orarr;':                           '↻'
	'&ord;':                             '⩝'
	'&#10845;':                          '⩝'
	'&order;':                           'ℴ'
	'&#8500;':                           'ℴ'
	'&orderof;':                         'ℴ'
	'&#170;':                            'ª'
	'&ordf;':                            'ª'
	'&#186;':                            'º'
	'&ordm;':                            'º'
	'&origof;':                          '⊶'
	'&#8886;':                           '⊶'
	'&oror;':                            '⩖'
	'&#10838;':                          '⩖'
	'&orslope;':                         '⩗'
	'&#10839;':                          '⩗'
	'&orv;':                             '⩛'
	'&#10843;':                          '⩛'
	'&oscr;':                            'ℴ'
	'&#248;':                            'ø'
	'&oslash;':                          'ø'
	'&osol;':                            '⊘'
	'&#8856;':                           '⊘'
	'&#245;':                            'õ'
	'&otilde;':                          'õ'
	'&otimes;':                          '⊗'
	'&otimesas;':                        '⨶'
	'&#10806;':                          '⨶'
	'&#246;':                            'ö'
	'&ouml;':                            'ö'
	'&ovbar;':                           '⌽'
	'&#9021;':                           '⌽'
	'&par;':                             '∥'
	'&#182;':                            '¶'
	'&para;':                            '¶'
	'&parallel;':                        '∥'
	'&parsim;':                          '⫳'
	'&#10995;':                          '⫳'
	'&parsl;':                           '⫽'
	'&#11005;':                          '⫽'
	'&part;':                            '∂'
	'&pcy;':                             'п'
	'&#1087;':                           'п'
	'&percnt;':                          '%'
	'&#37;':                             '%'
	'&period;':                          '.'
	'&#46;':                             '.'
	'&permil;':                          '‰'
	'&#8240;':                           '‰'
	'&perp;':                            '⊥'
	'&pertenk;':                         '‱'
	'&#8241;':                           '‱'
	'&pfr;':                             '𝔭'
	'&#120109;':                         '𝔭'
	'&phi;':                             'φ'
	'&#966;':                            'φ'
	'&phiv;':                            'ϕ'
	'&#981;':                            'ϕ'
	'&phmmat;':                          'ℳ'
	'&phone;':                           '☎'
	'&#9742;':                           '☎'
	'&pi;':                              'π'
	'&#960;':                            'π'
	'&pitchfork;':                       '⋔'
	'&piv;':                             'ϖ'
	'&#982;':                            'ϖ'
	'&planck;':                          'ℏ'
	'&planckh;':                         'ℎ'
	'&#8462;':                           'ℎ'
	'&plankv;':                          'ℏ'
	'&plus;':                            '+'
	'&#43;':                             '+'
	'&plusacir;':                        '⨣'
	'&#10787;':                          '⨣'
	'&plusb;':                           '⊞'
	'&pluscir;':                         '⨢'
	'&#10786;':                          '⨢'
	'&plusdo;':                          '∔'
	'&plusdu;':                          '⨥'
	'&#10789;':                          '⨥'
	'&pluse;':                           '⩲'
	'&#10866;':                          '⩲'
	'&plusmn;':                          '±'
	'&plussim;':                         '⨦'
	'&#10790;':                          '⨦'
	'&plustwo;':                         '⨧'
	'&#10791;':                          '⨧'
	'&pm;':                              '±'
	'&pointint;':                        '⨕'
	'&#10773;':                          '⨕'
	'&popf;':                            '𝕡'
	'&#120161;':                         '𝕡'
	'&#163;':                            '£'
	'&pound;':                           '£'
	'&pr;':                              '≺'
	'&prE;':                             '⪳'
	'&#10931;':                          '⪳'
	'&prap;':                            '⪷'
	'&#10935;':                          '⪷'
	'&prcue;':                           '≼'
	'&pre;':                             '⪯'
	'&prec;':                            '≺'
	'&precapprox;':                      '⪷'
	'&preccurlyeq;':                     '≼'
	'&preceq;':                          '⪯'
	'&precnapprox;':                     '⪹'
	'&#10937;':                          '⪹'
	'&precneqq;':                        '⪵'
	'&#10933;':                          '⪵'
	'&precnsim;':                        '⋨'
	'&#8936;':                           '⋨'
	'&precsim;':                         '≾'
	'&prime;':                           '′'
	'&#8242;':                           '′'
	'&primes;':                          'ℙ'
	'&prnE;':                            '⪵'
	'&prnap;':                           '⪹'
	'&prnsim;':                          '⋨'
	'&prod;':                            '∏'
	'&profalar;':                        '⌮'
	'&#9006;':                           '⌮'
	'&profline;':                        '⌒'
	'&#8978;':                           '⌒'
	'&profsurf;':                        '⌓'
	'&#8979;':                           '⌓'
	'&prop;':                            '∝'
	'&propto;':                          '∝'
	'&prsim;':                           '≾'
	'&prurel;':                          '⊰'
	'&#8880;':                           '⊰'
	'&pscr;':                            '𝓅'
	'&#120005;':                         '𝓅'
	'&psi;':                             'ψ'
	'&#968;':                            'ψ'
	'&puncsp;':                          ' '
	'&#8200;':                           ' '
	'&qfr;':                             '𝔮'
	'&#120110;':                         '𝔮'
	'&qint;':                            '⨌'
	'&qopf;':                            '𝕢'
	'&#120162;':                         '𝕢'
	'&qprime;':                          '⁗'
	'&#8279;':                           '⁗'
	'&qscr;':                            '𝓆'
	'&#120006;':                         '𝓆'
	'&quaternions;':                     'ℍ'
	'&quatint;':                         '⨖'
	'&#10774;':                          '⨖'
	'&quest;':                           '?'
	'&#63;':                             '?'
	'&questeq;':                         '≟'
	'&quot;':                            '"'
	'&rAarr;':                           '⇛'
	'&rArr;':                            '⇒'
	'&rAtail;':                          '⤜'
	'&#10524;':                          '⤜'
	'&rBarr;':                           '⤏'
	'&rHar;':                            '⥤'
	'&#10596;':                          '⥤'
	'&race;':                            '∽'
	'&#8765, 817;':                      '∽'
	'&racute;':                          'ŕ'
	'&#341;':                            'ŕ'
	'&radic;':                           '√'
	'&raemptyv;':                        '⦳'
	'&#10675;':                          '⦳'
	'&rang;':                            '⟩'
	'&rangd;':                           '⦒'
	'&#10642;':                          '⦒'
	'&range;':                           '⦥'
	'&#10661;':                          '⦥'
	'&rangle;':                          '⟩'
	'&#187;':                            '»'
	'&raquo;':                           '»'
	'&rarr;':                            '→'
	'&rarrap;':                          '⥵'
	'&#10613;':                          '⥵'
	'&rarrb;':                           '⇥'
	'&rarrbfs;':                         '⤠'
	'&#10528;':                          '⤠'
	'&rarrc;':                           '⤳'
	'&#10547;':                          '⤳'
	'&rarrfs;':                          '⤞'
	'&#10526;':                          '⤞'
	'&rarrhk;':                          '↪'
	'&rarrlp;':                          '↬'
	'&rarrpl;':                          '⥅'
	'&#10565;':                          '⥅'
	'&rarrsim;':                         '⥴'
	'&#10612;':                          '⥴'
	'&rarrtl;':                          '↣'
	'&#8611;':                           '↣'
	'&rarrw;':                           '↝'
	'&#8605;':                           '↝'
	'&ratail;':                          '⤚'
	'&#10522;':                          '⤚'
	'&ratio;':                           '∶'
	'&#8758;':                           '∶'
	'&rationals;':                       'ℚ'
	'&rbarr;':                           '⤍'
	'&rbbrk;':                           '❳'
	'&#10099;':                          '❳'
	'&rbrace;':                          '}'
	'&#125;':                            '}'
	'&rbrack;':                          ']'
	'&#93;':                             ']'
	'&rbrke;':                           '⦌'
	'&#10636;':                          '⦌'
	'&rbrksld;':                         '⦎'
	'&#10638;':                          '⦎'
	'&rbrkslu;':                         '⦐'
	'&#10640;':                          '⦐'
	'&rcaron;':                          'ř'
	'&#345;':                            'ř'
	'&rcedil;':                          'ŗ'
	'&#343;':                            'ŗ'
	'&rceil;':                           '⌉'
	'&rcub;':                            '}'
	'&rcy;':                             'р'
	'&#1088;':                           'р'
	'&rdca;':                            '⤷'
	'&#10551;':                          '⤷'
	'&rdldhar;':                         '⥩'
	'&#10601;':                          '⥩'
	'&rdquo;':                           '”'
	'&rdquor;':                          '”'
	'&rdsh;':                            '↳'
	'&#8627;':                           '↳'
	'&real;':                            'ℜ'
	'&realine;':                         'ℛ'
	'&realpart;':                        'ℜ'
	'&reals;':                           'ℝ'
	'&rect;':                            '▭'
	'&#9645;':                           '▭'
	'&reg;':                             '®'
	'&rfisht;':                          '⥽'
	'&#10621;':                          '⥽'
	'&rfloor;':                          '⌋'
	'&rfr;':                             '𝔯'
	'&#120111;':                         '𝔯'
	'&rhard;':                           '⇁'
	'&rharu;':                           '⇀'
	'&rharul;':                          '⥬'
	'&#10604;':                          '⥬'
	'&rho;':                             'ρ'
	'&#961;':                            'ρ'
	'&rhov;':                            'ϱ'
	'&#1009;':                           'ϱ'
	'&rightarrow;':                      '→'
	'&rightarrowtail;':                  '↣'
	'&rightharpoondown;':                '⇁'
	'&rightharpoonup;':                  '⇀'
	'&rightleftarrows;':                 '⇄'
	'&rightleftharpoons;':               '⇌'
	'&rightrightarrows;':                '⇉'
	'&#8649;':                           '⇉'
	'&rightsquigarrow;':                 '↝'
	'&rightthreetimes;':                 '⋌'
	'&#8908;':                           '⋌'
	'&ring;':                            '˚'
	'&#730;':                            '˚'
	'&risingdotseq;':                    '≓'
	'&rlarr;':                           '⇄'
	'&rlhar;':                           '⇌'
	'&rlm;':                             '‏'
	'&#8207;':                           '‏'
	'&rmoust;':                          '⎱'
	'&#9137;':                           '⎱'
	'&rmoustache;':                      '⎱'
	'&rnmid;':                           '⫮'
	'&#10990;':                          '⫮'
	'&roang;':                           '⟭'
	'&#10221;':                          '⟭'
	'&roarr;':                           '⇾'
	'&#8702;':                           '⇾'
	'&robrk;':                           '⟧'
	'&ropar;':                           '⦆'
	'&#10630;':                          '⦆'
	'&ropf;':                            '𝕣'
	'&#120163;':                         '𝕣'
	'&roplus;':                          '⨮'
	'&#10798;':                          '⨮'
	'&rotimes;':                         '⨵'
	'&#10805;':                          '⨵'
	'&rpar;':                            ')'
	'&#41;':                             ')'
	'&rpargt;':                          '⦔'
	'&#10644;':                          '⦔'
	'&rppolint;':                        '⨒'
	'&#10770;':                          '⨒'
	'&rrarr;':                           '⇉'
	'&rsaquo;':                          '›'
	'&#8250;':                           '›'
	'&rscr;':                            '𝓇'
	'&#120007;':                         '𝓇'
	'&rsh;':                             '↱'
	'&rsqb;':                            ']'
	'&rsquo;':                           '’'
	'&rsquor;':                          '’'
	'&rthree;':                          '⋌'
	'&rtimes;':                          '⋊'
	'&#8906;':                           '⋊'
	'&rtri;':                            '▹'
	'&#9657;':                           '▹'
	'&rtrie;':                           '⊵'
	'&rtrif;':                           '▸'
	'&rtriltri;':                        '⧎'
	'&#10702;':                          '⧎'
	'&ruluhar;':                         '⥨'
	'&#10600;':                          '⥨'
	'&rx;':                              '℞'
	'&#8478;':                           '℞'
	'&sacute;':                          'ś'
	'&#347;':                            'ś'
	'&sbquo;':                           '‚'
	'&sc;':                              '≻'
	'&scE;':                             '⪴'
	'&#10932;':                          '⪴'
	'&scap;':                            '⪸'
	'&#10936;':                          '⪸'
	'&scaron;':                          'š'
	'&#353;':                            'š'
	'&sccue;':                           '≽'
	'&sce;':                             '⪰'
	'&scedil;':                          'ş'
	'&#351;':                            'ş'
	'&scirc;':                           'ŝ'
	'&#349;':                            'ŝ'
	'&scnE;':                            '⪶'
	'&#10934;':                          '⪶'
	'&scnap;':                           '⪺'
	'&#10938;':                          '⪺'
	'&scnsim;':                          '⋩'
	'&#8937;':                           '⋩'
	'&scpolint;':                        '⨓'
	'&#10771;':                          '⨓'
	'&scsim;':                           '≿'
	'&scy;':                             'с'
	'&#1089;':                           'с'
	'&sdot;':                            '⋅'
	'&#8901;':                           '⋅'
	'&sdotb;':                           '⊡'
	'&sdote;':                           '⩦'
	'&#10854;':                          '⩦'
	'&seArr;':                           '⇘'
	'&#8664;':                           '⇘'
	'&searhk;':                          '⤥'
	'&searr;':                           '↘'
	'&searrow;':                         '↘'
	'&#167;':                            '§'
	'&sect;':                            '§'
	'&semi;':                            ';'
	'&#59;':                             ';'
	'&seswar;':                          '⤩'
	'&#10537;':                          '⤩'
	'&setminus;':                        '∖'
	'&setmn;':                           '∖'
	'&sext;':                            '✶'
	'&#10038;':                          '✶'
	'&sfr;':                             '𝔰'
	'&#120112;':                         '𝔰'
	'&sfrown;':                          '⌢'
	'&sharp;':                           '♯'
	'&#9839;':                           '♯'
	'&shchcy;':                          'щ'
	'&#1097;':                           'щ'
	'&shcy;':                            'ш'
	'&#1096;':                           'ш'
	'&shortmid;':                        '∣'
	'&shortparallel;':                   '∥'
	'&#173;':                            '­'
	'&shy;':                             '­'
	'&sigma;':                           'σ'
	'&#963;':                            'σ'
	'&sigmaf;':                          'ς'
	'&#962;':                            'ς'
	'&sigmav;':                          'ς'
	'&sim;':                             '∼'
	'&simdot;':                          '⩪'
	'&#10858;':                          '⩪'
	'&sime;':                            '≃'
	'&simeq;':                           '≃'
	'&simg;':                            '⪞'
	'&#10910;':                          '⪞'
	'&simgE;':                           '⪠'
	'&#10912;':                          '⪠'
	'&siml;':                            '⪝'
	'&#10909;':                          '⪝'
	'&simlE;':                           '⪟'
	'&#10911;':                          '⪟'
	'&simne;':                           '≆'
	'&#8774;':                           '≆'
	'&simplus;':                         '⨤'
	'&#10788;':                          '⨤'
	'&simrarr;':                         '⥲'
	'&#10610;':                          '⥲'
	'&slarr;':                           '←'
	'&smallsetminus;':                   '∖'
	'&smashp;':                          '⨳'
	'&#10803;':                          '⨳'
	'&smeparsl;':                        '⧤'
	'&#10724;':                          '⧤'
	'&smid;':                            '∣'
	'&smile;':                           '⌣'
	'&#8995;':                           '⌣'
	'&smt;':                             '⪪'
	'&#10922;':                          '⪪'
	'&smte;':                            '⪬'
	'&#10924;':                          '⪬'
	'&smtes;':                           '⪬'
	'&#10924, 65024;':                   '⪬'
	'&softcy;':                          'ь'
	'&#1100;':                           'ь'
	'&sol;':                             '/'
	'&#47;':                             '/'
	'&solb;':                            '⧄'
	'&#10692;':                          '⧄'
	'&solbar;':                          '⌿'
	'&#9023;':                           '⌿'
	'&sopf;':                            '𝕤'
	'&#120164;':                         '𝕤'
	'&spades;':                          '♠'
	'&#9824;':                           '♠'
	'&spadesuit;':                       '♠'
	'&spar;':                            '∥'
	'&sqcap;':                           '⊓'
	'&sqcaps;':                          '⊓'
	'&#8851, 65024;':                    '⊓'
	'&sqcup;':                           '⊔'
	'&sqcups;':                          '⊔'
	'&#8852, 65024;':                    '⊔'
	'&sqsub;':                           '⊏'
	'&sqsube;':                          '⊑'
	'&sqsubset;':                        '⊏'
	'&sqsubseteq;':                      '⊑'
	'&sqsup;':                           '⊐'
	'&sqsupe;':                          '⊒'
	'&sqsupset;':                        '⊐'
	'&sqsupseteq;':                      '⊒'
	'&squ;':                             '□'
	'&square;':                          '□'
	'&squarf;':                          '▪'
	'&squf;':                            '▪'
	'&srarr;':                           '→'
	'&sscr;':                            '𝓈'
	'&#120008;':                         '𝓈'
	'&ssetmn;':                          '∖'
	'&ssmile;':                          '⌣'
	'&sstarf;':                          '⋆'
	'&star;':                            '☆'
	'&#9734;':                           '☆'
	'&starf;':                           '★'
	'&straightepsilon;':                 'ϵ'
	'&straightphi;':                     'ϕ'
	'&strns;':                           '¯'
	'&sub;':                             '⊂'
	'&#8834;':                           '⊂'
	'&subE;':                            '⫅'
	'&#10949;':                          '⫅'
	'&subdot;':                          '⪽'
	'&#10941;':                          '⪽'
	'&sube;':                            '⊆'
	'&subedot;':                         '⫃'
	'&#10947;':                          '⫃'
	'&submult;':                         '⫁'
	'&#10945;':                          '⫁'
	'&subnE;':                           '⫋'
	'&#10955;':                          '⫋'
	'&subne;':                           '⊊'
	'&#8842;':                           '⊊'
	'&subplus;':                         '⪿'
	'&#10943;':                          '⪿'
	'&subrarr;':                         '⥹'
	'&#10617;':                          '⥹'
	'&subset;':                          '⊂'
	'&subseteq;':                        '⊆'
	'&subseteqq;':                       '⫅'
	'&subsetneq;':                       '⊊'
	'&subsetneqq;':                      '⫋'
	'&subsim;':                          '⫇'
	'&#10951;':                          '⫇'
	'&subsub;':                          '⫕'
	'&#10965;':                          '⫕'
	'&subsup;':                          '⫓'
	'&#10963;':                          '⫓'
	'&succ;':                            '≻'
	'&succapprox;':                      '⪸'
	'&succcurlyeq;':                     '≽'
	'&succeq;':                          '⪰'
	'&succnapprox;':                     '⪺'
	'&succneqq;':                        '⪶'
	'&succnsim;':                        '⋩'
	'&succsim;':                         '≿'
	'&sum;':                             '∑'
	'&sung;':                            '♪'
	'&#9834;':                           '♪'
	'&#185;':                            '¹'
	'&sup1;':                            '¹'
	'&#178;':                            '²'
	'&sup2;':                            '²'
	'&#179;':                            '³'
	'&sup3;':                            '³'
	'&sup;':                             '⊃'
	'&supE;':                            '⫆'
	'&#10950;':                          '⫆'
	'&supdot;':                          '⪾'
	'&#10942;':                          '⪾'
	'&supdsub;':                         '⫘'
	'&#10968;':                          '⫘'
	'&supe;':                            '⊇'
	'&supedot;':                         '⫄'
	'&#10948;':                          '⫄'
	'&suphsol;':                         '⟉'
	'&#10185;':                          '⟉'
	'&suphsub;':                         '⫗'
	'&#10967;':                          '⫗'
	'&suplarr;':                         '⥻'
	'&#10619;':                          '⥻'
	'&supmult;':                         '⫂'
	'&#10946;':                          '⫂'
	'&supnE;':                           '⫌'
	'&#10956;':                          '⫌'
	'&supne;':                           '⊋'
	'&#8843;':                           '⊋'
	'&supplus;':                         '⫀'
	'&#10944;':                          '⫀'
	'&supset;':                          '⊃'
	'&supseteq;':                        '⊇'
	'&supseteqq;':                       '⫆'
	'&supsetneq;':                       '⊋'
	'&supsetneqq;':                      '⫌'
	'&supsim;':                          '⫈'
	'&#10952;':                          '⫈'
	'&supsub;':                          '⫔'
	'&#10964;':                          '⫔'
	'&supsup;':                          '⫖'
	'&#10966;':                          '⫖'
	'&swArr;':                           '⇙'
	'&#8665;':                           '⇙'
	'&swarhk;':                          '⤦'
	'&swarr;':                           '↙'
	'&swarrow;':                         '↙'
	'&swnwar;':                          '⤪'
	'&#10538;':                          '⤪'
	'&#223;':                            'ß'
	'&szlig;':                           'ß'
	'&target;':                          '⌖'
	'&#8982;':                           '⌖'
	'&tau;':                             'τ'
	'&#964;':                            'τ'
	'&tbrk;':                            '⎴'
	'&tcaron;':                          'ť'
	'&#357;':                            'ť'
	'&tcedil;':                          'ţ'
	'&#355;':                            'ţ'
	'&tcy;':                             'т'
	'&#1090;':                           'т'
	'&tdot;':                            '⃛'
	'&telrec;':                          '⌕'
	'&#8981;':                           '⌕'
	'&tfr;':                             '𝔱'
	'&#120113;':                         '𝔱'
	'&there4;':                          '∴'
	'&therefore;':                       '∴'
	'&theta;':                           'θ'
	'&#952;':                            'θ'
	'&thetasym;':                        'ϑ'
	'&#977;':                            'ϑ'
	'&thetav;':                          'ϑ'
	'&thickapprox;':                     '≈'
	'&thicksim;':                        '∼'
	'&thinsp;':                          ' '
	'&thkap;':                           '≈'
	'&thksim;':                          '∼'
	'&#254;':                            'þ'
	'&thorn;':                           'þ'
	'&tilde;':                           '˜'
	'&#215;':                            '×'
	'&times;':                           '×'
	'&timesb;':                          '⊠'
	'&timesbar;':                        '⨱'
	'&#10801;':                          '⨱'
	'&timesd;':                          '⨰'
	'&#10800;':                          '⨰'
	'&tint;':                            '∭'
	'&toea;':                            '⤨'
	'&top;':                             '⊤'
	'&topbot;':                          '⌶'
	'&#9014;':                           '⌶'
	'&topcir;':                          '⫱'
	'&#10993;':                          '⫱'
	'&topf;':                            '𝕥'
	'&#120165;':                         '𝕥'
	'&topfork;':                         '⫚'
	'&#10970;':                          '⫚'
	'&tosa;':                            '⤩'
	'&tprime;':                          '‴'
	'&#8244;':                           '‴'
	'&trade;':                           '™'
	'&triangle;':                        '▵'
	'&#9653;':                           '▵'
	'&triangledown;':                    '▿'
	'&triangleleft;':                    '◃'
	'&trianglelefteq;':                  '⊴'
	'&triangleq;':                       '≜'
	'&#8796;':                           '≜'
	'&triangleright;':                   '▹'
	'&trianglerighteq;':                 '⊵'
	'&tridot;':                          '◬'
	'&#9708;':                           '◬'
	'&trie;':                            '≜'
	'&triminus;':                        '⨺'
	'&#10810;':                          '⨺'
	'&triplus;':                         '⨹'
	'&#10809;':                          '⨹'
	'&trisb;':                           '⧍'
	'&#10701;':                          '⧍'
	'&tritime;':                         '⨻'
	'&#10811;':                          '⨻'
	'&trpezium;':                        '⏢'
	'&#9186;':                           '⏢'
	'&tscr;':                            '𝓉'
	'&#120009;':                         '𝓉'
	'&tscy;':                            'ц'
	'&#1094;':                           'ц'
	'&tshcy;':                           'ћ'
	'&#1115;':                           'ћ'
	'&tstrok;':                          'ŧ'
	'&#359;':                            'ŧ'
	'&twixt;':                           '≬'
	'&twoheadleftarrow;':                '↞'
	'&twoheadrightarrow;':               '↠'
	'&uArr;':                            '⇑'
	'&uHar;':                            '⥣'
	'&#10595;':                          '⥣'
	'&#250;':                            'ú'
	'&uacute;':                          'ú'
	'&uarr;':                            '↑'
	'&ubrcy;':                           'ў'
	'&#1118;':                           'ў'
	'&ubreve;':                          'ŭ'
	'&#365;':                            'ŭ'
	'&#251;':                            'û'
	'&ucirc;':                           'û'
	'&ucy;':                             'у'
	'&#1091;':                           'у'
	'&udarr;':                           '⇅'
	'&udblac;':                          'ű'
	'&#369;':                            'ű'
	'&udhar;':                           '⥮'
	'&ufisht;':                          '⥾'
	'&#10622;':                          '⥾'
	'&ufr;':                             '𝔲'
	'&#120114;':                         '𝔲'
	'&#249;':                            'ù'
	'&ugrave;':                          'ù'
	'&uharl;':                           '↿'
	'&uharr;':                           '↾'
	'&uhblk;':                           '▀'
	'&#9600;':                           '▀'
	'&ulcorn;':                          '⌜'
	'&#8988;':                           '⌜'
	'&ulcorner;':                        '⌜'
	'&ulcrop;':                          '⌏'
	'&#8975;':                           '⌏'
	'&ultri;':                           '◸'
	'&#9720;':                           '◸'
	'&umacr;':                           'ū'
	'&#363;':                            'ū'
	'&uml;':                             '¨'
	'&uogon;':                           'ų'
	'&#371;':                            'ų'
	'&uopf;':                            '𝕦'
	'&#120166;':                         '𝕦'
	'&uparrow;':                         '↑'
	'&updownarrow;':                     '↕'
	'&upharpoonleft;':                   '↿'
	'&upharpoonright;':                  '↾'
	'&uplus;':                           '⊎'
	'&upsi;':                            'υ'
	'&#965;':                            'υ'
	'&upsih;':                           'ϒ'
	'&upsilon;':                         'υ'
	'&upuparrows;':                      '⇈'
	'&#8648;':                           '⇈'
	'&urcorn;':                          '⌝'
	'&#8989;':                           '⌝'
	'&urcorner;':                        '⌝'
	'&urcrop;':                          '⌎'
	'&#8974;':                           '⌎'
	'&uring;':                           'ů'
	'&#367;':                            'ů'
	'&urtri;':                           '◹'
	'&#9721;':                           '◹'
	'&uscr;':                            '𝓊'
	'&#120010;':                         '𝓊'
	'&utdot;':                           '⋰'
	'&#8944;':                           '⋰'
	'&utilde;':                          'ũ'
	'&#361;':                            'ũ'
	'&utri;':                            '▵'
	'&utrif;':                           '▴'
	'&uuarr;':                           '⇈'
	'&#252;':                            'ü'
	'&uuml;':                            'ü'
	'&uwangle;':                         '⦧'
	'&#10663;':                          '⦧'
	'&vArr;':                            '⇕'
	'&vBar;':                            '⫨'
	'&#10984;':                          '⫨'
	'&vBarv;':                           '⫩'
	'&#10985;':                          '⫩'
	'&vDash;':                           '⊨'
	'&vangrt;':                          '⦜'
	'&#10652;':                          '⦜'
	'&varepsilon;':                      'ϵ'
	'&varkappa;':                        'ϰ'
	'&varnothing;':                      '∅'
	'&varphi;':                          'ϕ'
	'&varpi;':                           'ϖ'
	'&varpropto;':                       '∝'
	'&varr;':                            '↕'
	'&varrho;':                          'ϱ'
	'&varsigma;':                        'ς'
	'&varsubsetneq;':                    '⊊'
	'&#8842, 65024;':                    '⊊'
	'&varsubsetneqq;':                   '⫋'
	'&#10955, 65024;':                   '⫋'
	'&varsupsetneq;':                    '⊋'
	'&#8843, 65024;':                    '⊋'
	'&varsupsetneqq;':                   '⫌'
	'&#10956, 65024;':                   '⫌'
	'&vartheta;':                        'ϑ'
	'&vartriangleleft;':                 '⊲'
	'&vartriangleright;':                '⊳'
	'&vcy;':                             'в'
	'&#1074;':                           'в'
	'&vdash;':                           '⊢'
	'&vee;':                             '∨'
	'&veebar;':                          '⊻'
	'&#8891;':                           '⊻'
	'&veeeq;':                           '≚'
	'&#8794;':                           '≚'
	'&vellip;':                          '⋮'
	'&#8942;':                           '⋮'
	'&verbar;':                          '|'
	'&vert;':                            '|'
	'&vfr;':                             '𝔳'
	'&#120115;':                         '𝔳'
	'&vltri;':                           '⊲'
	'&vnsub;':                           '⊂'
	'&vnsup;':                           '⊃'
	'&vopf;':                            '𝕧'
	'&#120167;':                         '𝕧'
	'&vprop;':                           '∝'
	'&vrtri;':                           '⊳'
	'&vscr;':                            '𝓋'
	'&#120011;':                         '𝓋'
	'&vsubnE;':                          '⫋'
	'&vsubne;':                          '⊊'
	'&vsupnE;':                          '⫌'
	'&vsupne;':                          '⊋'
	'&vzigzag;':                         '⦚'
	'&#10650;':                          '⦚'
	'&wcirc;':                           'ŵ'
	'&#373;':                            'ŵ'
	'&wedbar;':                          '⩟'
	'&#10847;':                          '⩟'
	'&wedge;':                           '∧'
	'&wedgeq;':                          '≙'
	'&#8793;':                           '≙'
	'&weierp;':                          '℘'
	'&#8472;':                           '℘'
	'&wfr;':                             '𝔴'
	'&#120116;':                         '𝔴'
	'&wopf;':                            '𝕨'
	'&#120168;':                         '𝕨'
	'&wp;':                              '℘'
	'&wr;':                              '≀'
	'&wreath;':                          '≀'
	'&wscr;':                            '𝓌'
	'&#120012;':                         '𝓌'
	'&xcap;':                            '⋂'
	'&xcirc;':                           '◯'
	'&xcup;':                            '⋃'
	'&xdtri;':                           '▽'
	'&xfr;':                             '𝔵'
	'&#120117;':                         '𝔵'
	'&xhArr;':                           '⟺'
	'&xharr;':                           '⟷'
	'&xi;':                              'ξ'
	'&#958;':                            'ξ'
	'&xlArr;':                           '⟸'
	'&xlarr;':                           '⟵'
	'&xmap;':                            '⟼'
	'&xnis;':                            '⋻'
	'&#8955;':                           '⋻'
	'&xodot;':                           '⨀'
	'&xopf;':                            '𝕩'
	'&#120169;':                         '𝕩'
	'&xoplus;':                          '⨁'
	'&xotime;':                          '⨂'
	'&xrArr;':                           '⟹'
	'&xrarr;':                           '⟶'
	'&xscr;':                            '𝓍'
	'&#120013;':                         '𝓍'
	'&xsqcup;':                          '⨆'
	'&xuplus;':                          '⨄'
	'&xutri;':                           '△'
	'&xvee;':                            '⋁'
	'&xwedge;':                          '⋀'
	'&#253;':                            'ý'
	'&yacute;':                          'ý'
	'&yacy;':                            'я'
	'&#1103;':                           'я'
	'&ycirc;':                           'ŷ'
	'&#375;':                            'ŷ'
	'&ycy;':                             'ы'
	'&#1099;':                           'ы'
	'&#165;':                            '¥'
	'&yen;':                             '¥'
	'&yfr;':                             '𝔶'
	'&#120118;':                         '𝔶'
	'&yicy;':                            'ї'
	'&#1111;':                           'ї'
	'&yopf;':                            '𝕪'
	'&#120170;':                         '𝕪'
	'&yscr;':                            '𝓎'
	'&#120014;':                         '𝓎'
	'&yucy;':                            'ю'
	'&#1102;':                           'ю'
	'&#255;':                            'ÿ'
	'&yuml;':                            'ÿ'
	'&zacute;':                          'ź'
	'&#378;':                            'ź'
	'&zcaron;':                          'ž'
	'&#382;':                            'ž'
	'&zcy;':                             'з'
	'&#1079;':                           'з'
	'&zdot;':                            'ż'
	'&#380;':                            'ż'
	'&zeetrf;':                          'ℨ'
	'&zeta;':                            'ζ'
	'&#950;':                            'ζ'
	'&zfr;':                             '𝔷'
	'&#120119;':                         '𝔷'
	'&zhcy;':                            'ж'
	'&#1078;':                           'ж'
	'&zigrarr;':                         '⇝'
	'&#8669;':                           '⇝'
	'&zopf;':                            '𝕫'
	'&#120171;':                         '𝕫'
	'&zscr;':                            '𝓏'
	'&#120015;':                         '𝓏'
	'&zwj;':                             '‍'
	'&#8205;':                           '‍'
	'&zwnj;':                            '‌'
	'&#8204;':                           '‌'
}

// htmlentity_to_string convert a html entity to its rune
pub fn htmlentity_to_string(data string) string {
	mut data_trasnform := data
	if data.contains('&') {
		for key, value in xmlreplacement.xml_replacement {
			data_trasnform = data_trasnform.replace(key, value)
		}
	}
	return data_transform
}
